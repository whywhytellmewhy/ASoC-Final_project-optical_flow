
//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_in_wait_coupled_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_coupled_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ../OpticalFlow_flow_calc.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Mon Jun 17 01:29:02 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, Flow_calc_COLUMN_C_14_tr0, Flow_calc_ROW_C_0_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [17:0] fsm_output;
  reg [17:0] fsm_output;
  input Flow_calc_COLUMN_C_14_tr0;
  input Flow_calc_ROW_C_0_tr0;


  // FSM State Type Declaration for OpticalFlow_flow_calc_run_run_fsm_1
  parameter
    main_C_0 = 5'd0,
    Flow_calc_COLUMN_C_0 = 5'd1,
    Flow_calc_COLUMN_C_1 = 5'd2,
    Flow_calc_COLUMN_C_2 = 5'd3,
    Flow_calc_COLUMN_C_3 = 5'd4,
    Flow_calc_COLUMN_C_4 = 5'd5,
    Flow_calc_COLUMN_C_5 = 5'd6,
    Flow_calc_COLUMN_C_6 = 5'd7,
    Flow_calc_COLUMN_C_7 = 5'd8,
    Flow_calc_COLUMN_C_8 = 5'd9,
    Flow_calc_COLUMN_C_9 = 5'd10,
    Flow_calc_COLUMN_C_10 = 5'd11,
    Flow_calc_COLUMN_C_11 = 5'd12,
    Flow_calc_COLUMN_C_12 = 5'd13,
    Flow_calc_COLUMN_C_13 = 5'd14,
    Flow_calc_COLUMN_C_14 = 5'd15,
    Flow_calc_ROW_C_0 = 5'd16,
    main_C_1 = 5'd17;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : OpticalFlow_flow_calc_run_run_fsm_1
    case (state_var)
      Flow_calc_COLUMN_C_0 : begin
        fsm_output = 18'b000000000000000010;
        state_var_NS = Flow_calc_COLUMN_C_1;
      end
      Flow_calc_COLUMN_C_1 : begin
        fsm_output = 18'b000000000000000100;
        state_var_NS = Flow_calc_COLUMN_C_2;
      end
      Flow_calc_COLUMN_C_2 : begin
        fsm_output = 18'b000000000000001000;
        state_var_NS = Flow_calc_COLUMN_C_3;
      end
      Flow_calc_COLUMN_C_3 : begin
        fsm_output = 18'b000000000000010000;
        state_var_NS = Flow_calc_COLUMN_C_4;
      end
      Flow_calc_COLUMN_C_4 : begin
        fsm_output = 18'b000000000000100000;
        state_var_NS = Flow_calc_COLUMN_C_5;
      end
      Flow_calc_COLUMN_C_5 : begin
        fsm_output = 18'b000000000001000000;
        state_var_NS = Flow_calc_COLUMN_C_6;
      end
      Flow_calc_COLUMN_C_6 : begin
        fsm_output = 18'b000000000010000000;
        state_var_NS = Flow_calc_COLUMN_C_7;
      end
      Flow_calc_COLUMN_C_7 : begin
        fsm_output = 18'b000000000100000000;
        state_var_NS = Flow_calc_COLUMN_C_8;
      end
      Flow_calc_COLUMN_C_8 : begin
        fsm_output = 18'b000000001000000000;
        state_var_NS = Flow_calc_COLUMN_C_9;
      end
      Flow_calc_COLUMN_C_9 : begin
        fsm_output = 18'b000000010000000000;
        state_var_NS = Flow_calc_COLUMN_C_10;
      end
      Flow_calc_COLUMN_C_10 : begin
        fsm_output = 18'b000000100000000000;
        state_var_NS = Flow_calc_COLUMN_C_11;
      end
      Flow_calc_COLUMN_C_11 : begin
        fsm_output = 18'b000001000000000000;
        state_var_NS = Flow_calc_COLUMN_C_12;
      end
      Flow_calc_COLUMN_C_12 : begin
        fsm_output = 18'b000010000000000000;
        state_var_NS = Flow_calc_COLUMN_C_13;
      end
      Flow_calc_COLUMN_C_13 : begin
        fsm_output = 18'b000100000000000000;
        state_var_NS = Flow_calc_COLUMN_C_14;
      end
      Flow_calc_COLUMN_C_14 : begin
        fsm_output = 18'b001000000000000000;
        if ( Flow_calc_COLUMN_C_14_tr0 ) begin
          state_var_NS = Flow_calc_ROW_C_0;
        end
        else begin
          state_var_NS = Flow_calc_COLUMN_C_0;
        end
      end
      Flow_calc_ROW_C_0 : begin
        fsm_output = 18'b010000000000000000;
        if ( Flow_calc_ROW_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = Flow_calc_COLUMN_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 18'b100000000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 18'b000000000000000001;
        state_var_NS = Flow_calc_COLUMN_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_run_staller
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_run_staller (
  run_wen, tensor_shift_rsci_wen_comp, shift_rsci_wen_comp, output_rsci_wen_comp
);
  output run_wen;
  input tensor_shift_rsci_wen_comp;
  input shift_rsci_wen_comp;
  input output_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = tensor_shift_rsci_wen_comp & shift_rsci_wen_comp & output_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_run_output_rsci_output_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_run_output_rsci_output_wait_ctrl (
  output_rsci_iswt0, output_rsci_biwt, output_rsci_irdy
);
  input output_rsci_iswt0;
  output output_rsci_biwt;
  input output_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_biwt = output_rsci_iswt0 & output_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_run_shift_rsci_shift_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_run_shift_rsci_shift_wait_ctrl (
  run_wen, shift_rsci_iswt0, shift_rsci_irdy_run_sct
);
  input run_wen;
  input shift_rsci_iswt0;
  output shift_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign shift_rsci_irdy_run_sct = shift_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_run_tensor_shift_rsci_tensor_shift_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_run_tensor_shift_rsci_tensor_shift_wait_ctrl (
  run_wen, tensor_shift_rsci_iswt0, tensor_shift_rsci_irdy_run_sct
);
  input run_wen;
  input tensor_shift_rsci_iswt0;
  output tensor_shift_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign tensor_shift_rsci_irdy_run_sct = tensor_shift_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_run_output_rsci
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_run_output_rsci (
  output_rsc_dat, output_rsc_vld, output_rsc_rdy, output_rsci_oswt, output_rsci_wen_comp,
      output_rsci_idat
);
  output [31:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input [31:0] output_rsci_idat;


  // Interconnect Declarations
  wire output_rsci_biwt;
  wire output_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd32)) output_rsci (
      .irdy(output_rsci_irdy),
      .ivld(output_rsci_oswt),
      .idat(output_rsci_idat),
      .rdy(output_rsc_rdy),
      .vld(output_rsc_vld),
      .dat(output_rsc_dat)
    );
  OpticalFlow_flow_calc_run_output_rsci_output_wait_ctrl OpticalFlow_flow_calc_run_output_rsci_output_wait_ctrl_inst
      (
      .output_rsci_iswt0(output_rsci_oswt),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_irdy(output_rsci_irdy)
    );
  assign output_rsci_wen_comp = (~ output_rsci_oswt) | output_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_run_shift_rsci
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_run_shift_rsci (
  shift_rsc_dat, shift_rsc_vld, shift_rsc_rdy, run_wen, shift_rsci_oswt, shift_rsci_wen_comp,
      shift_rsci_idat_mxwt
);
  input [8:0] shift_rsc_dat;
  input shift_rsc_vld;
  output shift_rsc_rdy;
  input run_wen;
  input shift_rsci_oswt;
  output shift_rsci_wen_comp;
  output [8:0] shift_rsci_idat_mxwt;


  // Interconnect Declarations
  wire shift_rsci_irdy_run_sct;
  wire shift_rsci_ivld;
  wire [8:0] shift_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd2),
  .width(32'sd9)) shift_rsci (
      .rdy(shift_rsc_rdy),
      .vld(shift_rsc_vld),
      .dat(shift_rsc_dat),
      .irdy(shift_rsci_irdy_run_sct),
      .ivld(shift_rsci_ivld),
      .idat(shift_rsci_idat)
    );
  OpticalFlow_flow_calc_run_shift_rsci_shift_wait_ctrl OpticalFlow_flow_calc_run_shift_rsci_shift_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .shift_rsci_iswt0(shift_rsci_oswt),
      .shift_rsci_irdy_run_sct(shift_rsci_irdy_run_sct)
    );
  assign shift_rsci_idat_mxwt = shift_rsci_idat;
  assign shift_rsci_wen_comp = (~ shift_rsci_oswt) | shift_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_run_tensor_shift_rsci
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_run_tensor_shift_rsci (
  tensor_shift_rsc_dat, tensor_shift_rsc_vld, tensor_shift_rsc_rdy, run_wen, tensor_shift_rsci_oswt,
      tensor_shift_rsci_wen_comp, tensor_shift_rsci_idat_mxwt
);
  input [191:0] tensor_shift_rsc_dat;
  input tensor_shift_rsc_vld;
  output tensor_shift_rsc_rdy;
  input run_wen;
  input tensor_shift_rsci_oswt;
  output tensor_shift_rsci_wen_comp;
  output [159:0] tensor_shift_rsci_idat_mxwt;


  // Interconnect Declarations
  wire tensor_shift_rsci_irdy_run_sct;
  wire tensor_shift_rsci_ivld;
  wire [191:0] tensor_shift_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd1),
  .width(32'sd192)) tensor_shift_rsci (
      .rdy(tensor_shift_rsc_rdy),
      .vld(tensor_shift_rsc_vld),
      .dat(tensor_shift_rsc_dat),
      .irdy(tensor_shift_rsci_irdy_run_sct),
      .ivld(tensor_shift_rsci_ivld),
      .idat(tensor_shift_rsci_idat)
    );
  OpticalFlow_flow_calc_run_tensor_shift_rsci_tensor_shift_wait_ctrl OpticalFlow_flow_calc_run_tensor_shift_rsci_tensor_shift_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .tensor_shift_rsci_iswt0(tensor_shift_rsci_oswt),
      .tensor_shift_rsci_irdy_run_sct(tensor_shift_rsci_irdy_run_sct)
    );
  assign tensor_shift_rsci_idat_mxwt = {(tensor_shift_rsci_idat[191:96]) , (tensor_shift_rsci_idat[63:0])};
  assign tensor_shift_rsci_wen_comp = (~ tensor_shift_rsci_oswt) | tensor_shift_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_run
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_run (
  clk, rst, arst_n, tensor_shift_rsc_dat, tensor_shift_rsc_vld, tensor_shift_rsc_rdy,
      shift_rsc_dat, shift_rsc_vld, shift_rsc_rdy, output_rsc_dat, output_rsc_vld,
      output_rsc_rdy, widthIn, heightIn, shift_threshold
);
  input clk;
  input rst;
  input arst_n;
  input [191:0] tensor_shift_rsc_dat;
  input tensor_shift_rsc_vld;
  output tensor_shift_rsc_rdy;
  input [8:0] shift_rsc_dat;
  input shift_rsc_vld;
  output shift_rsc_rdy;
  output [31:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  input [8:0] shift_threshold;


  // Interconnect Declarations
  wire run_wen;
  wire tensor_shift_rsci_wen_comp;
  wire [159:0] tensor_shift_rsci_idat_mxwt;
  wire shift_rsci_wen_comp;
  wire [8:0] shift_rsci_idat_mxwt;
  wire output_rsci_wen_comp;
  reg [31:0] output_rsci_idat;
  wire [17:0] fsm_output;
  wire Flow_calc_ROW_Flow_calc_ROW_if_Flow_calc_ROW_if_nor_tmp;
  wire Flow_calc_COLUMN_Flow_calc_COLUMN_if_1_Flow_calc_COLUMN_if_1_nor_tmp;
  wire or_dcpl_8;
  wire or_dcpl_10;
  wire or_dcpl_19;
  wire and_20_cse;
  wire and_21_cse;
  reg operator_9_false_slc_operator_9_false_acc_8_svs;
  reg Flow_calc_COLUMN_if_Flow_calc_COLUMN_if_and_2_itm;
  reg Flow_calc_COLUMN_if_if_slc_Flow_calc_COLUMN_if_if_acc_11_svs;
  wire tensor_shift_value_val_and_ssc;
  reg reg_output_rsci_iswt0_cse;
  reg reg_shift_rsci_iswt0_cse;
  wire Flow_calc_COLUMN_if_and_68_cse;
  wire Flow_calc_ROW_y_or_cse;
  wire [63:0] z_out;
  wire [63:0] z_out_1;
  reg [8:0] Flow_calc_ROW_y_sva;
  reg [10:0] Flow_calc_COLUMN_x_sva;
  reg [8:0] shift_value_sva;
  reg [63:0] denominator_value_sva;
  reg [63:0] velocity_value_x_sva;
  wire [64:0] nl_velocity_value_x_sva;
  reg [63:0] velocity_value_y_sva;
  wire [64:0] nl_velocity_value_y_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_28_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_26_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_25_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_35_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_24_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_36_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_22_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_19_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_16_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_44_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_45_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_46_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_12_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_48_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_10_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_50_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_52_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_54_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_56_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_58_sva;
  reg Flow_calc_COLUMN_if_and_2_psp_60_sva;
  reg [8:0] Flow_calc_COLUMN_if_ac_int_cctor_4_sva;
  reg [63:0] Flow_calc_COLUMN_if_sqr_itm;
  reg [63:0] Flow_calc_COLUMN_if_mul_2_itm;
  reg [63:0] Flow_calc_COLUMN_if_mul_3_itm;
  reg [63:0] Flow_calc_COLUMN_if_mul_4_itm;
  reg [4:0] operator_9_false_acc_44_itm;
  wire [5:0] nl_operator_9_false_acc_44_itm;
  reg [5:0] operator_9_false_acc_48_itm;
  wire [6:0] nl_operator_9_false_acc_48_itm;
  reg [8:0] operator_9_false_acc_83_itm;
  wire [12:0] nl_operator_9_false_acc_83_itm;
  reg [3:0] operator_9_false_acc_41_itm;
  wire [4:0] nl_operator_9_false_acc_41_itm;
  reg Flow_calc_COLUMN_if_and_57_itm;
  reg [2:0] operator_9_false_acc_39_itm;
  wire [3:0] nl_operator_9_false_acc_39_itm;
  reg Flow_calc_COLUMN_if_and_55_itm;
  reg Flow_calc_COLUMN_if_and_59_itm;
  reg Flow_calc_COLUMN_if_and_61_itm;
  reg [8:0] operator_9_false_acc_85_itm;
  wire [9:0] nl_operator_9_false_acc_85_itm;
  reg [8:0] operator_9_false_acc_84_itm;
  wire [11:0] nl_operator_9_false_acc_84_itm;
  reg [10:0] Flow_calc_COLUMN_acc_itm;
  wire [11:0] nl_Flow_calc_COLUMN_acc_itm;
  reg Flow_calc_COLUMN_if_and_2_seb;
  reg Flow_calc_COLUMN_if_and_3_seb;
  reg Flow_calc_COLUMN_if_and_7_seb;
  reg Flow_calc_COLUMN_if_and_33_seb;
  reg Flow_calc_COLUMN_if_and_49_seb;
  reg Flow_calc_COLUMN_if_and_seb;
  reg [1:0] operator_9_false_acc_94_cse;
  wire [2:0] nl_operator_9_false_acc_94_cse;
  reg [2:0] operator_9_false_acc_102_cse;
  wire [3:0] nl_operator_9_false_acc_102_cse;
  reg [3:0] operator_9_false_acc_57_itm_6_3;
  wire [4:0] nl_operator_9_false_acc_57_itm_6_3;
  reg [3:0] operator_9_false_acc_56_itm_6_3;
  wire [4:0] nl_operator_9_false_acc_56_itm_6_3;
  reg [4:0] operator_9_false_acc_55_itm_6_2;
  wire [5:0] nl_operator_9_false_acc_55_itm_6_2;
  reg [3:0] operator_9_false_acc_54_itm_6_3;
  wire [4:0] nl_operator_9_false_acc_54_itm_6_3;
  reg [4:0] operator_9_false_acc_53_itm_6_2;
  wire [5:0] nl_operator_9_false_acc_53_itm_6_2;
  reg [5:0] operator_9_false_acc_52_itm_6_1;
  wire [6:0] nl_operator_9_false_acc_52_itm_6_1;
  reg [3:0] operator_9_false_acc_45_itm_4_1;
  wire [4:0] nl_operator_9_false_acc_45_itm_4_1;
  reg [3:0] operator_9_false_acc_43_itm_4_1;
  wire [4:0] nl_operator_9_false_acc_43_itm_4_1;
  reg operator_9_false_acc_40_itm_1;
  reg [2:0] operator_9_false_acc_66_itm_2_0;
  wire [3:0] nl_operator_9_false_acc_66_itm_2_0;
  reg [5:0] operator_9_false_acc_65_itm_6_1;
  wire [6:0] nl_operator_9_false_acc_65_itm_6_1;
  reg [4:0] operator_9_false_acc_64_itm_6_2;
  wire [5:0] nl_operator_9_false_acc_64_itm_6_2;
  reg [3:0] operator_9_false_acc_63_itm_6_3;
  wire [4:0] nl_operator_9_false_acc_63_itm_6_3;
  reg [1:0] operator_9_false_acc_63_itm_2_1;
  wire [2:0] nl_operator_9_false_acc_63_itm_2_1;
  reg [3:0] operator_9_false_acc_62_itm_6_3;
  wire [4:0] nl_operator_9_false_acc_62_itm_6_3;
  reg [2:0] operator_9_false_acc_60_itm_6_4;
  wire [3:0] nl_operator_9_false_acc_60_itm_6_4;
  reg [1:0] operator_9_false_acc_60_itm_3_2;
  wire [2:0] nl_operator_9_false_acc_60_itm_3_2;
  reg [2:0] operator_9_false_acc_59_itm_6_4;
  wire [3:0] nl_operator_9_false_acc_59_itm_6_4;
  reg [1:0] operator_9_false_acc_59_itm_2_1;
  wire [2:0] nl_operator_9_false_acc_59_itm_2_1;
  reg [2:0] operator_9_false_acc_58_itm_6_4;
  wire [3:0] nl_operator_9_false_acc_58_itm_6_4;
  wire output_rsci_idat_mx0c0;
  wire Flow_calc_COLUMN_if_and_2_psp_48_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_50_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_52_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_54_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_56_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_58_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_60_sva_1;
  wire Flow_calc_COLUMN_if_and_seb_1;
  wire Flow_calc_COLUMN_if_and_49_seb_1;
  wire Flow_calc_COLUMN_if_and_2_psp_19_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_10_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_22_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_44_sva_1;
  wire Flow_calc_COLUMN_if_and_33_seb_1;
  wire Flow_calc_COLUMN_if_and_2_psp_45_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_12_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_16_sva_1;
  wire Flow_calc_COLUMN_if_and_7_seb_1;
  wire Flow_calc_COLUMN_if_and_2_psp_26_sva_1;
  wire Flow_calc_COLUMN_if_and_3_seb_1;
  wire Flow_calc_COLUMN_if_and_2_psp_35_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_28_sva_1;
  wire Flow_calc_COLUMN_if_and_2_seb_1;
  wire Flow_calc_COLUMN_if_and_2_psp_25_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_24_sva_1;
  wire [63:0] denominator_value_sva_1;
  wire [64:0] nl_denominator_value_sva_1;
  wire Flow_calc_COLUMN_if_for_16_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire [62:0] Flow_calc_COLUMN_if_acc_6_sdt_sva_1;
  wire [63:0] nl_Flow_calc_COLUMN_if_acc_6_sdt_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_49_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_51_sva_1;
  wire Flow_calc_COLUMN_if_for_10_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_8_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_57_sva_1;
  wire Flow_calc_COLUMN_if_for_4_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_2_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_1_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_41_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_32_sva_1;
  wire Flow_calc_COLUMN_if_for_63_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_62_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_60_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_9_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_4_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_17_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_8_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_33_sva_1;
  wire Flow_calc_COLUMN_if_for_61_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_39_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_42_sva_1;
  wire Flow_calc_COLUMN_if_for_58_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_57_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_34_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_20_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_21_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_43_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_18_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_38_sva_1;
  wire Flow_calc_COLUMN_if_for_56_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_and_2_psp_37_sva_1;
  wire Flow_calc_COLUMN_if_for_50_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_49_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_48_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_52_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_36_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_34_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_40_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_33_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire velocity_value_compare_to_sign_bit_bitwise_OR_complement_35_32_sva_1;
  wire Flow_calc_COLUMN_if_for_3_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_5_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_6_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_7_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_59_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_9_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_11_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_55_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_12_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_54_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_13_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_53_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_14_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_15_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_51_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_17_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_18_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_19_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_47_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_20_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_46_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_21_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_45_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_22_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_44_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_23_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_43_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_24_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_42_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_25_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_41_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_26_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_27_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_39_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_28_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_38_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_29_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_37_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire Flow_calc_COLUMN_if_for_30_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire velocity_value_compare_to_sign_bit_bitwise_OR_complement_35_33_sva_1;
  wire Flow_calc_COLUMN_if_for_35_Flow_calc_COLUMN_if_for_or_1_psp_sva_1;
  wire operator_9_false_asn_76;
  wire [8:0] Flow_calc_COLUMN_if_ac_int_cctor_4_sva_1;
  wire [9:0] nl_Flow_calc_COLUMN_if_ac_int_cctor_4_sva_1;
  wire [9:0] Flow_calc_COLUMN_if_if_acc_1_sdt_1;
  wire [10:0] nl_Flow_calc_COLUMN_if_if_acc_1_sdt_1;
  wire [11:0] operator_11_false_1_acc_psp_sva_1;
  wire [12:0] nl_operator_11_false_1_acc_psp_sva_1;
  wire [9:0] operator_9_false_2_acc_psp_sva_1;
  wire [10:0] nl_operator_9_false_2_acc_psp_sva_1;
  reg [95:0] tensor_shift_value_val_sva_191_96;
  reg [63:0] tensor_shift_value_val_sva_63_0;
  wire operator_11_false_acc_itm_12_1;
  wire operator_11_false_acc_itm_10_1;
  wire operator_9_false_acc_itm_10_1;

  wire[31:0] Flow_calc_COLUMN_if_if_nand_nl;
  wire Flow_calc_COLUMN_if_if_not_9_nl;
  wire Flow_calc_COLUMN_x_not_1_nl;
  wire[8:0] Flow_calc_ROW_acc_nl;
  wire[9:0] nl_Flow_calc_ROW_acc_nl;
  wire Flow_calc_ROW_y_not_1_nl;
  wire[8:0] operator_9_false_acc_nl;
  wire[9:0] nl_operator_9_false_acc_nl;
  wire Flow_calc_COLUMN_if_and_36_nl;
  wire Flow_calc_COLUMN_if_and_48_nl;
  wire Flow_calc_COLUMN_if_and_52_nl;
  wire Flow_calc_COLUMN_if_and_60_nl;
  wire Flow_calc_COLUMN_if_and_1_nl;
  wire Flow_calc_COLUMN_if_and_51_nl;
  wire Flow_calc_COLUMN_if_and_47_nl;
  wire Flow_calc_COLUMN_if_and_35_nl;
  wire Flow_calc_COLUMN_if_and_31_nl;
  wire Flow_calc_COLUMN_if_and_39_nl;
  wire Flow_calc_COLUMN_if_and_15_nl;
  wire Flow_calc_COLUMN_if_and_4_nl;
  wire[3:0] operator_9_false_acc_109_nl;
  wire[4:0] nl_operator_9_false_acc_109_nl;
  wire[2:0] operator_9_false_acc_110_nl;
  wire[3:0] nl_operator_9_false_acc_110_nl;
  wire[8:0] operator_9_false_acc_82_nl;
  wire[9:0] nl_operator_9_false_acc_82_nl;
  wire[6:0] operator_9_false_acc_51_nl;
  wire[8:0] nl_operator_9_false_acc_51_nl;
  wire[6:0] operator_9_false_acc_69_nl;
  wire[7:0] nl_operator_9_false_acc_69_nl;
  wire[4:0] operator_9_false_acc_49_nl;
  wire[5:0] nl_operator_9_false_acc_49_nl;
  wire[7:0] operator_9_false_acc_77_nl;
  wire[10:0] nl_operator_9_false_acc_77_nl;
  wire[11:0] Flow_calc_COLUMN_if_if_acc_nl;
  wire[12:0] nl_Flow_calc_COLUMN_if_if_acc_nl;
  wire[9:0] Flow_calc_COLUMN_if_if_acc_3_nl;
  wire[10:0] nl_Flow_calc_COLUMN_if_if_acc_3_nl;
  wire[12:0] operator_11_false_acc_nl;
  wire[13:0] nl_operator_11_false_acc_nl;
  wire[11:0] operator_11_false_acc_1_nl;
  wire[12:0] nl_operator_11_false_acc_1_nl;
  wire[10:0] operator_11_false_acc_nl_1;
  wire[11:0] nl_operator_11_false_acc_nl_1;
  wire[10:0] operator_9_false_acc_nl_1;
  wire[11:0] nl_operator_9_false_acc_nl_1;
  wire[9:0] operator_9_false_acc_1_nl;
  wire[10:0] nl_operator_9_false_acc_1_nl;
  wire[8:0] operator_9_false_acc_nl_2;
  wire[9:0] nl_operator_9_false_acc_nl_2;
  wire[31:0] Flow_calc_COLUMN_if_mux1h_39_nl;
  wire Flow_calc_COLUMN_if_or_5_nl;
  wire Flow_calc_COLUMN_if_or_6_nl;
  wire[31:0] Flow_calc_COLUMN_if_mux1h_40_nl;
  wire Flow_calc_COLUMN_if_or_7_nl;
  wire Flow_calc_COLUMN_if_or_8_nl;
  wire signed [63:0] nl_mul_sgnd;

  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_Flow_calc_COLUMN_if_lshift_rg_a;
  assign nl_Flow_calc_COLUMN_if_lshift_rg_a = MUX1HOT_v_64_3_2(denominator_value_sva,
      velocity_value_x_sva, velocity_value_y_sva, {(fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14])});
  mgc_shift_l_v5 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd64)) Flow_calc_COLUMN_if_lshift_rg (
      .a(nl_Flow_calc_COLUMN_if_lshift_rg_a[63:0]),
      .s(Flow_calc_COLUMN_if_ac_int_cctor_4_sva),
      .z(z_out)
    );
  OpticalFlow_flow_calc_run_tensor_shift_rsci OpticalFlow_flow_calc_run_tensor_shift_rsci_inst
      (
      .tensor_shift_rsc_dat(tensor_shift_rsc_dat),
      .tensor_shift_rsc_vld(tensor_shift_rsc_vld),
      .tensor_shift_rsc_rdy(tensor_shift_rsc_rdy),
      .run_wen(run_wen),
      .tensor_shift_rsci_oswt(reg_shift_rsci_iswt0_cse),
      .tensor_shift_rsci_wen_comp(tensor_shift_rsci_wen_comp),
      .tensor_shift_rsci_idat_mxwt(tensor_shift_rsci_idat_mxwt)
    );
  OpticalFlow_flow_calc_run_shift_rsci OpticalFlow_flow_calc_run_shift_rsci_inst
      (
      .shift_rsc_dat(shift_rsc_dat),
      .shift_rsc_vld(shift_rsc_vld),
      .shift_rsc_rdy(shift_rsc_rdy),
      .run_wen(run_wen),
      .shift_rsci_oswt(reg_shift_rsci_iswt0_cse),
      .shift_rsci_wen_comp(shift_rsci_wen_comp),
      .shift_rsci_idat_mxwt(shift_rsci_idat_mxwt)
    );
  OpticalFlow_flow_calc_run_output_rsci OpticalFlow_flow_calc_run_output_rsci_inst
      (
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .output_rsci_oswt(reg_output_rsci_iswt0_cse),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_idat(output_rsci_idat)
    );
  OpticalFlow_flow_calc_run_staller OpticalFlow_flow_calc_run_staller_inst (
      .run_wen(run_wen),
      .tensor_shift_rsci_wen_comp(tensor_shift_rsci_wen_comp),
      .shift_rsci_wen_comp(shift_rsci_wen_comp),
      .output_rsci_wen_comp(output_rsci_wen_comp)
    );
  OpticalFlow_flow_calc_run_run_fsm OpticalFlow_flow_calc_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .Flow_calc_COLUMN_C_14_tr0(Flow_calc_COLUMN_Flow_calc_COLUMN_if_1_Flow_calc_COLUMN_if_1_nor_tmp),
      .Flow_calc_ROW_C_0_tr0(Flow_calc_ROW_Flow_calc_ROW_if_Flow_calc_ROW_if_nor_tmp)
    );
  assign Flow_calc_ROW_y_or_cse = (fsm_output[0]) | (fsm_output[16]);
  assign tensor_shift_value_val_and_ssc = run_wen & (~(or_dcpl_10 | (fsm_output[3])
      | or_dcpl_8 | (fsm_output[6])));
  assign Flow_calc_COLUMN_if_and_68_cse = run_wen & (fsm_output[13:12]==2'b00);
  assign nl_operator_11_false_acc_1_nl = conv_u2u_11_12(Flow_calc_COLUMN_x_sva) +
      conv_u2u_11_12(~ widthIn);
  assign operator_11_false_acc_1_nl = nl_operator_11_false_acc_1_nl[11:0];
  assign nl_operator_11_false_acc_nl = conv_u2s_12_13(operator_11_false_acc_1_nl)
      + 13'b1100000000011;
  assign operator_11_false_acc_nl = nl_operator_11_false_acc_nl[12:0];
  assign operator_11_false_acc_itm_12_1 = readslicef_13_1_12(operator_11_false_acc_nl);
  assign nl_operator_11_false_acc_nl_1 = conv_u2u_10_11(Flow_calc_COLUMN_x_sva[10:1])
      + 11'b11111111111;
  assign operator_11_false_acc_nl_1 = nl_operator_11_false_acc_nl_1[10:0];
  assign operator_11_false_acc_itm_10_1 = readslicef_11_1_10(operator_11_false_acc_nl_1);
  assign nl_operator_9_false_acc_1_nl = conv_u2u_9_10(Flow_calc_ROW_y_sva) + conv_u2u_9_10(~
      heightIn);
  assign operator_9_false_acc_1_nl = nl_operator_9_false_acc_1_nl[9:0];
  assign nl_operator_9_false_acc_nl_1 = conv_u2s_10_11(operator_9_false_acc_1_nl)
      + 11'b11000000011;
  assign operator_9_false_acc_nl_1 = nl_operator_9_false_acc_nl_1[10:0];
  assign operator_9_false_acc_itm_10_1 = readslicef_11_1_10(operator_9_false_acc_nl_1);
  assign Flow_calc_COLUMN_if_and_2_psp_48_sva_1 = Flow_calc_COLUMN_if_for_15_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[48]);
  assign Flow_calc_COLUMN_if_and_2_psp_50_sva_1 = Flow_calc_COLUMN_if_for_13_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[50]);
  assign Flow_calc_COLUMN_if_and_2_psp_52_sva_1 = Flow_calc_COLUMN_if_for_11_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[52]);
  assign Flow_calc_COLUMN_if_and_2_psp_54_sva_1 = Flow_calc_COLUMN_if_for_9_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[54]);
  assign Flow_calc_COLUMN_if_and_2_psp_56_sva_1 = Flow_calc_COLUMN_if_for_7_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[56]);
  assign Flow_calc_COLUMN_if_and_2_psp_58_sva_1 = Flow_calc_COLUMN_if_for_5_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[58]);
  assign Flow_calc_COLUMN_if_and_2_psp_60_sva_1 = Flow_calc_COLUMN_if_for_3_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[60]);
  assign Flow_calc_COLUMN_if_and_seb_1 = Flow_calc_COLUMN_if_for_1_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[62]);
  assign Flow_calc_COLUMN_if_and_49_seb_1 = Flow_calc_COLUMN_if_for_57_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[6]);
  assign Flow_calc_COLUMN_if_and_2_psp_19_sva_1 = Flow_calc_COLUMN_if_for_44_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[19]);
  assign Flow_calc_COLUMN_if_and_2_psp_10_sva_1 = Flow_calc_COLUMN_if_for_53_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[10]);
  assign Flow_calc_COLUMN_if_and_2_psp_22_sva_1 = Flow_calc_COLUMN_if_for_41_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[22]);
  assign Flow_calc_COLUMN_if_and_2_psp_44_sva_1 = Flow_calc_COLUMN_if_for_19_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[44]);
  assign Flow_calc_COLUMN_if_and_33_seb_1 = Flow_calc_COLUMN_if_for_49_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[14]);
  assign Flow_calc_COLUMN_if_and_2_psp_45_sva_1 = Flow_calc_COLUMN_if_for_18_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[45]);
  assign Flow_calc_COLUMN_if_and_2_psp_12_sva_1 = Flow_calc_COLUMN_if_for_51_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[12]);
  assign Flow_calc_COLUMN_if_and_2_psp_16_sva_1 = Flow_calc_COLUMN_if_for_47_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[16]);
  assign Flow_calc_COLUMN_if_and_7_seb_1 = Flow_calc_COLUMN_if_for_36_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[27]);
  assign Flow_calc_COLUMN_if_and_2_psp_26_sva_1 = Flow_calc_COLUMN_if_for_37_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[26]);
  assign Flow_calc_COLUMN_if_and_3_seb_1 = Flow_calc_COLUMN_if_for_34_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[29]);
  assign Flow_calc_COLUMN_if_and_2_psp_35_sva_1 = Flow_calc_COLUMN_if_for_28_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[35]);
  assign Flow_calc_COLUMN_if_and_2_psp_28_sva_1 = Flow_calc_COLUMN_if_for_35_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[28]);
  assign Flow_calc_COLUMN_if_and_2_seb_1 = Flow_calc_COLUMN_if_for_33_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[30]);
  assign Flow_calc_COLUMN_if_and_2_psp_25_sva_1 = Flow_calc_COLUMN_if_for_38_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[25]);
  assign Flow_calc_COLUMN_if_and_2_psp_24_sva_1 = Flow_calc_COLUMN_if_for_39_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[24]);
  assign nl_denominator_value_sva_1 = Flow_calc_COLUMN_if_mul_3_itm - Flow_calc_COLUMN_if_sqr_itm;
  assign denominator_value_sva_1 = nl_denominator_value_sva_1[63:0];
  assign Flow_calc_COLUMN_if_for_16_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[15])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[15]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[15]));
  assign nl_Flow_calc_COLUMN_if_acc_6_sdt_sva_1 = ({(~ Flow_calc_COLUMN_if_for_1_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_2_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_3_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_4_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_5_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_6_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_7_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_8_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_9_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_10_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_11_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_12_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_13_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_14_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_15_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_16_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_17_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_18_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_19_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_20_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_21_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_22_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_23_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_24_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_25_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_26_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_27_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_28_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_29_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_30_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ velocity_value_compare_to_sign_bit_bitwise_OR_complement_35_33_sva_1)
      , (~ velocity_value_compare_to_sign_bit_bitwise_OR_complement_35_32_sva_1)
      , (~ Flow_calc_COLUMN_if_for_33_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_34_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_35_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_36_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_37_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_38_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_39_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_40_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_41_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_42_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_43_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_44_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_45_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_46_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_47_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_48_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_49_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_50_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_51_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_52_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_53_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_54_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_55_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_56_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_57_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_58_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_59_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_60_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~
      Flow_calc_COLUMN_if_for_61_Flow_calc_COLUMN_if_for_or_1_psp_sva_1) , (~ Flow_calc_COLUMN_if_for_62_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)
      , (~ Flow_calc_COLUMN_if_for_63_Flow_calc_COLUMN_if_for_or_1_psp_sva_1)}) +
      63'b000000000000000000000000000000000000000000000000000000000000001;
  assign Flow_calc_COLUMN_if_acc_6_sdt_sva_1 = nl_Flow_calc_COLUMN_if_acc_6_sdt_sva_1[62:0];
  assign Flow_calc_COLUMN_if_and_2_psp_49_sva_1 = Flow_calc_COLUMN_if_for_14_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[49]);
  assign Flow_calc_COLUMN_if_and_2_psp_51_sva_1 = Flow_calc_COLUMN_if_for_12_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[51]);
  assign Flow_calc_COLUMN_if_for_10_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[9])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[9]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[9]));
  assign Flow_calc_COLUMN_if_for_8_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[7])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[7]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[7]));
  assign Flow_calc_COLUMN_if_and_2_psp_57_sva_1 = Flow_calc_COLUMN_if_for_6_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[57]);
  assign Flow_calc_COLUMN_if_for_4_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[3])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[3]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[3]));
  assign Flow_calc_COLUMN_if_for_2_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[1])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[1]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[1]));
  assign Flow_calc_COLUMN_if_for_1_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[0])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[0]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[0]));
  assign Flow_calc_COLUMN_if_and_2_psp_41_sva_1 = Flow_calc_COLUMN_if_for_22_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[41]);
  assign Flow_calc_COLUMN_if_and_2_psp_32_sva_1 = velocity_value_compare_to_sign_bit_bitwise_OR_complement_35_33_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[32]);
  assign Flow_calc_COLUMN_if_for_63_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[62])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[62]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[62]));
  assign Flow_calc_COLUMN_if_for_62_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[61])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[61]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[61]));
  assign Flow_calc_COLUMN_if_for_60_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[59])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[59]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[59]));
  assign Flow_calc_COLUMN_if_and_2_psp_9_sva_1 = Flow_calc_COLUMN_if_for_54_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[9]);
  assign Flow_calc_COLUMN_if_and_2_psp_4_sva_1 = Flow_calc_COLUMN_if_for_59_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[4]);
  assign Flow_calc_COLUMN_if_and_2_psp_17_sva_1 = Flow_calc_COLUMN_if_for_46_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[17]);
  assign Flow_calc_COLUMN_if_and_2_psp_8_sva_1 = Flow_calc_COLUMN_if_for_55_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[8]);
  assign Flow_calc_COLUMN_if_and_2_psp_33_sva_1 = Flow_calc_COLUMN_if_for_30_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[33]);
  assign Flow_calc_COLUMN_if_for_61_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[60])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[60]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[60]));
  assign Flow_calc_COLUMN_if_and_2_psp_39_sva_1 = Flow_calc_COLUMN_if_for_24_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[39]);
  assign Flow_calc_COLUMN_if_and_2_psp_42_sva_1 = Flow_calc_COLUMN_if_for_21_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[42]);
  assign Flow_calc_COLUMN_if_for_58_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[57])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[57]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[57]));
  assign Flow_calc_COLUMN_if_for_57_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[56])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[56]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[56]));
  assign Flow_calc_COLUMN_if_and_2_psp_34_sva_1 = Flow_calc_COLUMN_if_for_29_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[34]);
  assign Flow_calc_COLUMN_if_and_2_psp_20_sva_1 = Flow_calc_COLUMN_if_for_43_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[20]);
  assign Flow_calc_COLUMN_if_and_2_psp_21_sva_1 = Flow_calc_COLUMN_if_for_42_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[21]);
  assign Flow_calc_COLUMN_if_and_2_psp_43_sva_1 = Flow_calc_COLUMN_if_for_20_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[43]);
  assign Flow_calc_COLUMN_if_and_2_psp_18_sva_1 = Flow_calc_COLUMN_if_for_45_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[18]);
  assign Flow_calc_COLUMN_if_and_2_psp_38_sva_1 = Flow_calc_COLUMN_if_for_25_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[38]);
  assign Flow_calc_COLUMN_if_for_56_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[55])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[55]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[55]));
  assign Flow_calc_COLUMN_if_and_2_psp_37_sva_1 = Flow_calc_COLUMN_if_for_26_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[37]);
  assign Flow_calc_COLUMN_if_for_50_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[49])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[49]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[49]));
  assign Flow_calc_COLUMN_if_for_49_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[48])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[48]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[48]));
  assign Flow_calc_COLUMN_if_for_48_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[47])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[47]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[47]));
  assign Flow_calc_COLUMN_if_for_52_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[51])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[51]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[51]));
  assign Flow_calc_COLUMN_if_for_36_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[35])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[35]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[35]));
  assign Flow_calc_COLUMN_if_for_34_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[33])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[33]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[33]));
  assign Flow_calc_COLUMN_if_for_40_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[39])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[39]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[39]));
  assign Flow_calc_COLUMN_if_for_33_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[32])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[32]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[32]));
  assign velocity_value_compare_to_sign_bit_bitwise_OR_complement_35_32_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[31])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[31]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[31]));
  assign Flow_calc_COLUMN_if_for_3_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[2])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[2]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[2]));
  assign Flow_calc_COLUMN_if_for_5_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[4])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[4]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[4]));
  assign Flow_calc_COLUMN_if_for_6_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[5])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[5]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[5]));
  assign Flow_calc_COLUMN_if_for_7_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[6])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[6]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[6]));
  assign Flow_calc_COLUMN_if_for_59_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[58])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[58]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[58]));
  assign Flow_calc_COLUMN_if_for_9_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[8])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[8]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[8]));
  assign Flow_calc_COLUMN_if_for_11_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[10])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[10]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[10]));
  assign Flow_calc_COLUMN_if_for_55_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[54])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[54]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[54]));
  assign Flow_calc_COLUMN_if_for_12_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[11])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[11]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[11]));
  assign Flow_calc_COLUMN_if_for_54_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[53])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[53]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[53]));
  assign Flow_calc_COLUMN_if_for_13_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[12])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[12]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[12]));
  assign Flow_calc_COLUMN_if_for_53_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[52])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[52]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[52]));
  assign Flow_calc_COLUMN_if_for_14_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[13])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[13]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[13]));
  assign Flow_calc_COLUMN_if_for_15_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[14])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[14]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[14]));
  assign Flow_calc_COLUMN_if_for_51_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[50])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[50]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[50]));
  assign Flow_calc_COLUMN_if_for_17_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[16])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[16]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[16]));
  assign Flow_calc_COLUMN_if_for_18_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[17])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[17]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[17]));
  assign Flow_calc_COLUMN_if_for_19_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[18])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[18]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[18]));
  assign Flow_calc_COLUMN_if_for_47_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[46])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[46]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[46]));
  assign Flow_calc_COLUMN_if_for_20_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[19])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[19]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[19]));
  assign Flow_calc_COLUMN_if_for_46_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[45])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[45]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[45]));
  assign Flow_calc_COLUMN_if_for_21_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[20])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[20]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[20]));
  assign Flow_calc_COLUMN_if_for_45_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[44])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[44]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[44]));
  assign Flow_calc_COLUMN_if_for_22_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[21])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[21]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[21]));
  assign Flow_calc_COLUMN_if_for_44_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[43])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[43]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[43]));
  assign Flow_calc_COLUMN_if_for_23_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[22])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[22]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[22]));
  assign Flow_calc_COLUMN_if_for_43_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[42])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[42]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[42]));
  assign Flow_calc_COLUMN_if_for_24_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[23])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[23]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[23]));
  assign Flow_calc_COLUMN_if_for_42_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[41])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[41]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[41]));
  assign Flow_calc_COLUMN_if_for_25_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[24])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[24]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[24]));
  assign Flow_calc_COLUMN_if_for_41_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[40])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[40]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[40]));
  assign Flow_calc_COLUMN_if_for_26_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[25])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[25]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[25]));
  assign Flow_calc_COLUMN_if_for_27_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[26])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[26]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[26]));
  assign Flow_calc_COLUMN_if_for_39_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[38])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[38]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[38]));
  assign Flow_calc_COLUMN_if_for_28_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[27])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[27]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[27]));
  assign Flow_calc_COLUMN_if_for_38_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[37])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[37]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[37]));
  assign Flow_calc_COLUMN_if_for_29_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[28])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[28]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[28]));
  assign Flow_calc_COLUMN_if_for_37_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[36])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[36]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[36]));
  assign Flow_calc_COLUMN_if_for_30_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[29])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[29]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[29]));
  assign velocity_value_compare_to_sign_bit_bitwise_OR_complement_35_33_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[30])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[30]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[30]));
  assign Flow_calc_COLUMN_if_for_35_Flow_calc_COLUMN_if_for_or_1_psp_sva_1 = ((denominator_value_sva_1[63])
      ^ (denominator_value_sva_1[34])) | ((velocity_value_x_sva[63]) ^ (velocity_value_x_sva[34]))
      | ((velocity_value_y_sva[63]) ^ (velocity_value_y_sva[34]));
  assign operator_9_false_asn_76 = Flow_calc_COLUMN_if_for_23_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[40]);
  assign nl_operator_9_false_acc_nl_2 = operator_9_false_acc_83_itm + operator_9_false_acc_85_itm;
  assign operator_9_false_acc_nl_2 = nl_operator_9_false_acc_nl_2[8:0];
  assign nl_Flow_calc_COLUMN_if_ac_int_cctor_4_sva_1 = operator_9_false_acc_nl_2
      + operator_9_false_acc_84_itm;
  assign Flow_calc_COLUMN_if_ac_int_cctor_4_sva_1 = nl_Flow_calc_COLUMN_if_ac_int_cctor_4_sva_1[8:0];
  assign nl_Flow_calc_COLUMN_if_if_acc_1_sdt_1 = conv_u2u_9_10(shift_threshold) +
      conv_u2u_9_10(~ Flow_calc_COLUMN_if_ac_int_cctor_4_sva_1);
  assign Flow_calc_COLUMN_if_if_acc_1_sdt_1 = nl_Flow_calc_COLUMN_if_if_acc_1_sdt_1[9:0];
  assign nl_operator_11_false_1_acc_psp_sva_1 = conv_u2s_11_12(widthIn) + 12'b111111111111;
  assign operator_11_false_1_acc_psp_sva_1 = nl_operator_11_false_1_acc_psp_sva_1[11:0];
  assign nl_operator_9_false_2_acc_psp_sva_1 = conv_u2s_9_10(heightIn) + 10'b1111111111;
  assign operator_9_false_2_acc_psp_sva_1 = nl_operator_9_false_2_acc_psp_sva_1[9:0];
  assign Flow_calc_ROW_Flow_calc_ROW_if_Flow_calc_ROW_if_nor_tmp = ~((Flow_calc_ROW_y_sva
      != (operator_9_false_2_acc_psp_sva_1[8:0])) | (operator_9_false_2_acc_psp_sva_1[9]));
  assign Flow_calc_COLUMN_Flow_calc_COLUMN_if_1_Flow_calc_COLUMN_if_1_nor_tmp = ~((Flow_calc_COLUMN_x_sva
      != (operator_11_false_1_acc_psp_sva_1[10:0])) | (operator_11_false_1_acc_psp_sva_1[11]));
  assign or_dcpl_8 = (fsm_output[2]) | (fsm_output[4]);
  assign or_dcpl_10 = (fsm_output[5]) | (fsm_output[7]);
  assign or_dcpl_19 = (fsm_output[8]) | (fsm_output[12]);
  assign and_20_cse = ~(Flow_calc_COLUMN_if_Flow_calc_COLUMN_if_and_2_itm | (~((fsm_output[4:3]!=2'b00))));
  assign and_21_cse = ((~ operator_9_false_acc_itm_10_1) | operator_9_false_slc_operator_9_false_acc_8_svs
      | (~((~ operator_11_false_acc_itm_10_1) & operator_11_false_acc_itm_12_1)))
      & (fsm_output[2]);
  assign output_rsci_idat_mx0c0 = and_20_cse | and_21_cse;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      output_rsci_idat <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      output_rsci_idat <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & (output_rsci_idat_mx0c0 | (Flow_calc_COLUMN_if_Flow_calc_COLUMN_if_and_2_itm
        & (fsm_output[12])) | (Flow_calc_COLUMN_if_Flow_calc_COLUMN_if_and_2_itm
        & (fsm_output[13])) | (Flow_calc_COLUMN_if_Flow_calc_COLUMN_if_and_2_itm
        & (fsm_output[14]))) ) begin
      output_rsci_idat <= ~(MUX_v_32_2_2(Flow_calc_COLUMN_if_if_nand_nl, 32'b11111111111111111111111111111111,
          output_rsci_idat_mx0c0));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Flow_calc_COLUMN_x_sva <= 11'b00000000000;
    end
    else if ( rst ) begin
      Flow_calc_COLUMN_x_sva <= 11'b00000000000;
    end
    else if ( run_wen & ((fsm_output[15]) | Flow_calc_ROW_y_or_cse) ) begin
      Flow_calc_COLUMN_x_sva <= MUX_v_11_2_2(11'b00000000000, Flow_calc_COLUMN_acc_itm,
          Flow_calc_COLUMN_x_not_1_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Flow_calc_ROW_y_sva <= 9'b000000000;
    end
    else if ( rst ) begin
      Flow_calc_ROW_y_sva <= 9'b000000000;
    end
    else if ( run_wen & Flow_calc_ROW_y_or_cse ) begin
      Flow_calc_ROW_y_sva <= MUX_v_9_2_2(9'b000000000, Flow_calc_ROW_acc_nl, Flow_calc_ROW_y_not_1_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_output_rsci_iswt0_cse <= 1'b0;
      reg_shift_rsci_iswt0_cse <= 1'b0;
      operator_9_false_slc_operator_9_false_acc_8_svs <= 1'b0;
      Flow_calc_COLUMN_if_mul_3_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      operator_9_false_acc_58_itm_6_4 <= 3'b000;
      Flow_calc_COLUMN_if_and_2_psp_48_sva <= 1'b0;
      operator_9_false_acc_59_itm_6_4 <= 3'b000;
      Flow_calc_COLUMN_if_and_2_psp_50_sva <= 1'b0;
      operator_9_false_acc_59_itm_2_1 <= 2'b00;
      operator_9_false_acc_60_itm_6_4 <= 3'b000;
      Flow_calc_COLUMN_if_and_2_psp_52_sva <= 1'b0;
      operator_9_false_acc_60_itm_3_2 <= 2'b00;
      operator_9_false_acc_102_cse <= 3'b000;
      Flow_calc_COLUMN_if_and_2_psp_54_sva <= 1'b0;
      operator_9_false_acc_62_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_psp_56_sva <= 1'b0;
      operator_9_false_acc_63_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_psp_58_sva <= 1'b0;
      operator_9_false_acc_63_itm_2_1 <= 2'b00;
      operator_9_false_acc_64_itm_6_2 <= 5'b00000;
      Flow_calc_COLUMN_if_and_2_psp_60_sva <= 1'b0;
      operator_9_false_acc_65_itm_6_1 <= 6'b000000;
      Flow_calc_COLUMN_if_and_seb <= 1'b0;
      operator_9_false_acc_66_itm_2_0 <= 3'b000;
      operator_9_false_acc_94_cse <= 2'b00;
      Flow_calc_COLUMN_if_and_61_itm <= 1'b0;
      Flow_calc_COLUMN_if_and_59_itm <= 1'b0;
      Flow_calc_COLUMN_if_and_55_itm <= 1'b0;
      operator_9_false_acc_39_itm <= 3'b000;
      operator_9_false_acc_40_itm_1 <= 1'b0;
      Flow_calc_COLUMN_if_and_57_itm <= 1'b0;
      operator_9_false_acc_43_itm_4_1 <= 4'b0000;
      Flow_calc_COLUMN_if_and_49_seb <= 1'b0;
      operator_9_false_acc_41_itm <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_psp_19_sva <= 1'b0;
      operator_9_false_acc_48_itm <= 6'b000000;
      operator_9_false_acc_44_itm <= 5'b00000;
      Flow_calc_COLUMN_if_and_2_psp_10_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_22_sva <= 1'b0;
      operator_9_false_acc_45_itm_4_1 <= 4'b0000;
      operator_9_false_acc_52_itm_6_1 <= 6'b000000;
      Flow_calc_COLUMN_if_and_2_psp_44_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_33_seb <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_45_sva <= 1'b0;
      operator_9_false_acc_53_itm_6_2 <= 5'b00000;
      Flow_calc_COLUMN_if_and_2_psp_12_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_16_sva <= 1'b0;
      operator_9_false_acc_54_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_7_seb <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_26_sva <= 1'b0;
      operator_9_false_acc_55_itm_6_2 <= 5'b00000;
      Flow_calc_COLUMN_if_and_3_seb <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_35_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_28_sva <= 1'b0;
      operator_9_false_acc_56_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_seb <= 1'b0;
      operator_9_false_acc_57_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_psp_25_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_24_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_46_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_36_sva <= 1'b0;
      operator_9_false_acc_84_itm <= 9'b000000000;
      operator_9_false_acc_85_itm <= 9'b000000000;
      operator_9_false_acc_83_itm <= 9'b000000000;
    end
    else if ( rst ) begin
      reg_output_rsci_iswt0_cse <= 1'b0;
      reg_shift_rsci_iswt0_cse <= 1'b0;
      operator_9_false_slc_operator_9_false_acc_8_svs <= 1'b0;
      Flow_calc_COLUMN_if_mul_3_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      operator_9_false_acc_58_itm_6_4 <= 3'b000;
      Flow_calc_COLUMN_if_and_2_psp_48_sva <= 1'b0;
      operator_9_false_acc_59_itm_6_4 <= 3'b000;
      Flow_calc_COLUMN_if_and_2_psp_50_sva <= 1'b0;
      operator_9_false_acc_59_itm_2_1 <= 2'b00;
      operator_9_false_acc_60_itm_6_4 <= 3'b000;
      Flow_calc_COLUMN_if_and_2_psp_52_sva <= 1'b0;
      operator_9_false_acc_60_itm_3_2 <= 2'b00;
      operator_9_false_acc_102_cse <= 3'b000;
      Flow_calc_COLUMN_if_and_2_psp_54_sva <= 1'b0;
      operator_9_false_acc_62_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_psp_56_sva <= 1'b0;
      operator_9_false_acc_63_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_psp_58_sva <= 1'b0;
      operator_9_false_acc_63_itm_2_1 <= 2'b00;
      operator_9_false_acc_64_itm_6_2 <= 5'b00000;
      Flow_calc_COLUMN_if_and_2_psp_60_sva <= 1'b0;
      operator_9_false_acc_65_itm_6_1 <= 6'b000000;
      Flow_calc_COLUMN_if_and_seb <= 1'b0;
      operator_9_false_acc_66_itm_2_0 <= 3'b000;
      operator_9_false_acc_94_cse <= 2'b00;
      Flow_calc_COLUMN_if_and_61_itm <= 1'b0;
      Flow_calc_COLUMN_if_and_59_itm <= 1'b0;
      Flow_calc_COLUMN_if_and_55_itm <= 1'b0;
      operator_9_false_acc_39_itm <= 3'b000;
      operator_9_false_acc_40_itm_1 <= 1'b0;
      Flow_calc_COLUMN_if_and_57_itm <= 1'b0;
      operator_9_false_acc_43_itm_4_1 <= 4'b0000;
      Flow_calc_COLUMN_if_and_49_seb <= 1'b0;
      operator_9_false_acc_41_itm <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_psp_19_sva <= 1'b0;
      operator_9_false_acc_48_itm <= 6'b000000;
      operator_9_false_acc_44_itm <= 5'b00000;
      Flow_calc_COLUMN_if_and_2_psp_10_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_22_sva <= 1'b0;
      operator_9_false_acc_45_itm_4_1 <= 4'b0000;
      operator_9_false_acc_52_itm_6_1 <= 6'b000000;
      Flow_calc_COLUMN_if_and_2_psp_44_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_33_seb <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_45_sva <= 1'b0;
      operator_9_false_acc_53_itm_6_2 <= 5'b00000;
      Flow_calc_COLUMN_if_and_2_psp_12_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_16_sva <= 1'b0;
      operator_9_false_acc_54_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_7_seb <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_26_sva <= 1'b0;
      operator_9_false_acc_55_itm_6_2 <= 5'b00000;
      Flow_calc_COLUMN_if_and_3_seb <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_35_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_28_sva <= 1'b0;
      operator_9_false_acc_56_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_seb <= 1'b0;
      operator_9_false_acc_57_itm_6_3 <= 4'b0000;
      Flow_calc_COLUMN_if_and_2_psp_25_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_24_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_46_sva <= 1'b0;
      Flow_calc_COLUMN_if_and_2_psp_36_sva <= 1'b0;
      operator_9_false_acc_84_itm <= 9'b000000000;
      operator_9_false_acc_85_itm <= 9'b000000000;
      operator_9_false_acc_83_itm <= 9'b000000000;
    end
    else if ( run_wen ) begin
      reg_output_rsci_iswt0_cse <= and_20_cse | (Flow_calc_COLUMN_if_Flow_calc_COLUMN_if_and_2_itm
          & ((fsm_output[14:12]!=3'b000))) | and_21_cse;
      reg_shift_rsci_iswt0_cse <= ~((Flow_calc_COLUMN_Flow_calc_COLUMN_if_1_Flow_calc_COLUMN_if_1_nor_tmp
          & (fsm_output[15])) | (~((fsm_output[15]) | (fsm_output[0]) | (fsm_output[16])))
          | (Flow_calc_ROW_Flow_calc_ROW_if_Flow_calc_ROW_if_nor_tmp & (fsm_output[16])));
      operator_9_false_slc_operator_9_false_acc_8_svs <= readslicef_9_1_8(operator_9_false_acc_nl);
      Flow_calc_COLUMN_if_mul_3_itm <= z_out_1;
      operator_9_false_acc_58_itm_6_4 <= nl_operator_9_false_acc_58_itm_6_4[2:0];
      Flow_calc_COLUMN_if_and_2_psp_48_sva <= Flow_calc_COLUMN_if_and_2_psp_48_sva_1;
      operator_9_false_acc_59_itm_6_4 <= nl_operator_9_false_acc_59_itm_6_4[2:0];
      Flow_calc_COLUMN_if_and_2_psp_50_sva <= Flow_calc_COLUMN_if_and_2_psp_50_sva_1;
      operator_9_false_acc_59_itm_2_1 <= nl_operator_9_false_acc_59_itm_2_1[1:0];
      operator_9_false_acc_60_itm_6_4 <= nl_operator_9_false_acc_60_itm_6_4[2:0];
      Flow_calc_COLUMN_if_and_2_psp_52_sva <= Flow_calc_COLUMN_if_and_2_psp_52_sva_1;
      operator_9_false_acc_60_itm_3_2 <= nl_operator_9_false_acc_60_itm_3_2[1:0];
      operator_9_false_acc_102_cse <= nl_operator_9_false_acc_102_cse[2:0];
      Flow_calc_COLUMN_if_and_2_psp_54_sva <= Flow_calc_COLUMN_if_and_2_psp_54_sva_1;
      operator_9_false_acc_62_itm_6_3 <= nl_operator_9_false_acc_62_itm_6_3[3:0];
      Flow_calc_COLUMN_if_and_2_psp_56_sva <= Flow_calc_COLUMN_if_and_2_psp_56_sva_1;
      operator_9_false_acc_63_itm_6_3 <= nl_operator_9_false_acc_63_itm_6_3[3:0];
      Flow_calc_COLUMN_if_and_2_psp_58_sva <= Flow_calc_COLUMN_if_and_2_psp_58_sva_1;
      operator_9_false_acc_63_itm_2_1 <= nl_operator_9_false_acc_63_itm_2_1[1:0];
      operator_9_false_acc_64_itm_6_2 <= nl_operator_9_false_acc_64_itm_6_2[4:0];
      Flow_calc_COLUMN_if_and_2_psp_60_sva <= Flow_calc_COLUMN_if_and_2_psp_60_sva_1;
      operator_9_false_acc_65_itm_6_1 <= nl_operator_9_false_acc_65_itm_6_1[5:0];
      Flow_calc_COLUMN_if_and_seb <= Flow_calc_COLUMN_if_and_seb_1;
      operator_9_false_acc_66_itm_2_0 <= nl_operator_9_false_acc_66_itm_2_0[2:0];
      operator_9_false_acc_94_cse <= nl_operator_9_false_acc_94_cse[1:0];
      Flow_calc_COLUMN_if_and_61_itm <= Flow_calc_COLUMN_if_for_63_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
          & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[0]);
      Flow_calc_COLUMN_if_and_59_itm <= Flow_calc_COLUMN_if_for_62_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
          & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[1]);
      Flow_calc_COLUMN_if_and_55_itm <= Flow_calc_COLUMN_if_for_60_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
          & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[3]);
      operator_9_false_acc_39_itm <= nl_operator_9_false_acc_39_itm[2:0];
      operator_9_false_acc_40_itm_1 <= ~ Flow_calc_COLUMN_if_and_2_psp_33_sva_1;
      Flow_calc_COLUMN_if_and_57_itm <= Flow_calc_COLUMN_if_for_61_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
          & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[2]);
      operator_9_false_acc_43_itm_4_1 <= nl_operator_9_false_acc_43_itm_4_1[3:0];
      Flow_calc_COLUMN_if_and_49_seb <= Flow_calc_COLUMN_if_and_49_seb_1;
      operator_9_false_acc_41_itm <= nl_operator_9_false_acc_41_itm[3:0];
      Flow_calc_COLUMN_if_and_2_psp_19_sva <= Flow_calc_COLUMN_if_and_2_psp_19_sva_1;
      operator_9_false_acc_48_itm <= nl_operator_9_false_acc_48_itm[5:0];
      operator_9_false_acc_44_itm <= nl_operator_9_false_acc_44_itm[4:0];
      Flow_calc_COLUMN_if_and_2_psp_10_sva <= Flow_calc_COLUMN_if_and_2_psp_10_sva_1;
      Flow_calc_COLUMN_if_and_2_psp_22_sva <= Flow_calc_COLUMN_if_and_2_psp_22_sva_1;
      operator_9_false_acc_45_itm_4_1 <= nl_operator_9_false_acc_45_itm_4_1[3:0];
      operator_9_false_acc_52_itm_6_1 <= nl_operator_9_false_acc_52_itm_6_1[5:0];
      Flow_calc_COLUMN_if_and_2_psp_44_sva <= Flow_calc_COLUMN_if_and_2_psp_44_sva_1;
      Flow_calc_COLUMN_if_and_33_seb <= Flow_calc_COLUMN_if_and_33_seb_1;
      Flow_calc_COLUMN_if_and_2_psp_45_sva <= Flow_calc_COLUMN_if_and_2_psp_45_sva_1;
      operator_9_false_acc_53_itm_6_2 <= nl_operator_9_false_acc_53_itm_6_2[4:0];
      Flow_calc_COLUMN_if_and_2_psp_12_sva <= Flow_calc_COLUMN_if_and_2_psp_12_sva_1;
      Flow_calc_COLUMN_if_and_2_psp_16_sva <= Flow_calc_COLUMN_if_and_2_psp_16_sva_1;
      operator_9_false_acc_54_itm_6_3 <= nl_operator_9_false_acc_54_itm_6_3[3:0];
      Flow_calc_COLUMN_if_and_7_seb <= Flow_calc_COLUMN_if_and_7_seb_1;
      Flow_calc_COLUMN_if_and_2_psp_26_sva <= Flow_calc_COLUMN_if_and_2_psp_26_sva_1;
      operator_9_false_acc_55_itm_6_2 <= nl_operator_9_false_acc_55_itm_6_2[4:0];
      Flow_calc_COLUMN_if_and_3_seb <= Flow_calc_COLUMN_if_and_3_seb_1;
      Flow_calc_COLUMN_if_and_2_psp_35_sva <= Flow_calc_COLUMN_if_and_2_psp_35_sva_1;
      Flow_calc_COLUMN_if_and_2_psp_28_sva <= Flow_calc_COLUMN_if_and_2_psp_28_sva_1;
      operator_9_false_acc_56_itm_6_3 <= nl_operator_9_false_acc_56_itm_6_3[3:0];
      Flow_calc_COLUMN_if_and_2_seb <= Flow_calc_COLUMN_if_and_2_seb_1;
      operator_9_false_acc_57_itm_6_3 <= nl_operator_9_false_acc_57_itm_6_3[3:0];
      Flow_calc_COLUMN_if_and_2_psp_25_sva <= Flow_calc_COLUMN_if_and_2_psp_25_sva_1;
      Flow_calc_COLUMN_if_and_2_psp_24_sva <= Flow_calc_COLUMN_if_and_2_psp_24_sva_1;
      Flow_calc_COLUMN_if_and_2_psp_46_sva <= Flow_calc_COLUMN_if_for_17_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
          & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[46]);
      Flow_calc_COLUMN_if_and_2_psp_36_sva <= Flow_calc_COLUMN_if_for_27_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
          & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[36]);
      operator_9_false_acc_84_itm <= nl_operator_9_false_acc_84_itm[8:0];
      operator_9_false_acc_85_itm <= nl_operator_9_false_acc_85_itm[8:0];
      operator_9_false_acc_83_itm <= nl_operator_9_false_acc_83_itm[8:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      tensor_shift_value_val_sva_191_96 <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      tensor_shift_value_val_sva_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      tensor_shift_value_val_sva_191_96 <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      tensor_shift_value_val_sva_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( tensor_shift_value_val_and_ssc ) begin
      tensor_shift_value_val_sva_191_96 <= tensor_shift_rsci_idat_mxwt[159:64];
      tensor_shift_value_val_sva_63_0 <= tensor_shift_rsci_idat_mxwt[63:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      shift_value_sva <= 9'b000000000;
    end
    else if ( rst ) begin
      shift_value_sva <= 9'b000000000;
    end
    else if ( run_wen & (~(or_dcpl_10 | (fsm_output[9]) | (fsm_output[10]) | (fsm_output[3])
        | or_dcpl_8 | (fsm_output[6]) | (fsm_output[8]))) ) begin
      shift_value_sva <= shift_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Flow_calc_COLUMN_acc_itm <= 11'b00000000000;
    end
    else if ( rst ) begin
      Flow_calc_COLUMN_acc_itm <= 11'b00000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      Flow_calc_COLUMN_acc_itm <= nl_Flow_calc_COLUMN_acc_itm[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Flow_calc_COLUMN_if_Flow_calc_COLUMN_if_and_2_itm <= 1'b0;
    end
    else if ( rst ) begin
      Flow_calc_COLUMN_if_Flow_calc_COLUMN_if_and_2_itm <= 1'b0;
    end
    else if ( run_wen & (fsm_output[2]) ) begin
      Flow_calc_COLUMN_if_Flow_calc_COLUMN_if_and_2_itm <= operator_11_false_acc_itm_12_1
          & (~ operator_11_false_acc_itm_10_1) & operator_9_false_acc_itm_10_1 &
          (~ operator_9_false_slc_operator_9_false_acc_8_svs);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Flow_calc_COLUMN_if_mul_4_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      Flow_calc_COLUMN_if_mul_4_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~ (fsm_output[4])) ) begin
      Flow_calc_COLUMN_if_mul_4_itm <= z_out_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      velocity_value_y_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      velocity_value_y_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((fsm_output[7]) | (fsm_output[11]) | (fsm_output[9]) |
        (fsm_output[10]) | (fsm_output[13]) | (fsm_output[6]) | or_dcpl_19)) ) begin
      velocity_value_y_sva <= nl_velocity_value_y_sva[63:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Flow_calc_COLUMN_if_mul_2_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      Flow_calc_COLUMN_if_mul_2_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~ (fsm_output[6])) ) begin
      Flow_calc_COLUMN_if_mul_2_itm <= z_out_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      velocity_value_x_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      velocity_value_x_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((fsm_output[11:9]!=3'b000) | or_dcpl_19)) ) begin
      velocity_value_x_sva <= nl_velocity_value_x_sva[63:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Flow_calc_COLUMN_if_sqr_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      Flow_calc_COLUMN_if_sqr_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~ (fsm_output[8])) ) begin
      Flow_calc_COLUMN_if_sqr_itm <= z_out_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      denominator_value_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      denominator_value_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[11:10]==2'b00) ) begin
      denominator_value_sva <= denominator_value_sva_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Flow_calc_COLUMN_if_ac_int_cctor_4_sva <= 9'b000000000;
      Flow_calc_COLUMN_if_if_slc_Flow_calc_COLUMN_if_if_acc_11_svs <= 1'b0;
    end
    else if ( rst ) begin
      Flow_calc_COLUMN_if_ac_int_cctor_4_sva <= 9'b000000000;
      Flow_calc_COLUMN_if_if_slc_Flow_calc_COLUMN_if_if_acc_11_svs <= 1'b0;
    end
    else if ( Flow_calc_COLUMN_if_and_68_cse ) begin
      Flow_calc_COLUMN_if_ac_int_cctor_4_sva <= Flow_calc_COLUMN_if_ac_int_cctor_4_sva_1;
      Flow_calc_COLUMN_if_if_slc_Flow_calc_COLUMN_if_if_acc_11_svs <= readslicef_12_1_11(Flow_calc_COLUMN_if_if_acc_nl);
    end
  end
  assign Flow_calc_COLUMN_if_if_not_9_nl = ~ Flow_calc_COLUMN_if_if_slc_Flow_calc_COLUMN_if_if_acc_11_svs;
  assign Flow_calc_COLUMN_if_if_nand_nl = ~(MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (z_out[63:32]), Flow_calc_COLUMN_if_if_not_9_nl));
  assign Flow_calc_COLUMN_x_not_1_nl = ~ Flow_calc_ROW_y_or_cse;
  assign nl_Flow_calc_ROW_acc_nl = Flow_calc_ROW_y_sva + 9'b000000001;
  assign Flow_calc_ROW_acc_nl = nl_Flow_calc_ROW_acc_nl[8:0];
  assign Flow_calc_ROW_y_not_1_nl = ~ (fsm_output[0]);
  assign nl_operator_9_false_acc_nl = conv_u2u_8_9(Flow_calc_ROW_y_sva[8:1]) + 9'b111111111;
  assign operator_9_false_acc_nl = nl_operator_9_false_acc_nl[8:0];
  assign Flow_calc_COLUMN_if_and_36_nl = Flow_calc_COLUMN_if_for_16_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[47]);
  assign nl_operator_9_false_acc_58_itm_6_4  = conv_u2u_2_3({{1{Flow_calc_COLUMN_if_and_2_psp_48_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_48_sva_1}) + conv_u2u_2_3(signext_2_1(Flow_calc_COLUMN_if_and_36_nl));
  assign nl_operator_9_false_acc_59_itm_6_4  = conv_u2u_2_3({{1{Flow_calc_COLUMN_if_and_2_psp_50_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_50_sva_1}) + conv_u2u_2_3({{1{Flow_calc_COLUMN_if_and_2_psp_49_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_49_sva_1});
  assign nl_operator_9_false_acc_59_itm_2_1  = conv_u2u_1_2(Flow_calc_COLUMN_if_and_2_psp_50_sva_1)
      + conv_u2u_1_2(Flow_calc_COLUMN_if_and_2_psp_49_sva_1);
  assign nl_operator_9_false_acc_60_itm_6_4  = conv_u2u_2_3({{1{Flow_calc_COLUMN_if_and_2_psp_52_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_52_sva_1}) + conv_u2u_2_3({{1{Flow_calc_COLUMN_if_and_2_psp_51_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_51_sva_1});
  assign nl_operator_9_false_acc_60_itm_3_2  = conv_u2u_1_2(Flow_calc_COLUMN_if_and_2_psp_52_sva_1)
      + conv_u2u_1_2(Flow_calc_COLUMN_if_and_2_psp_51_sva_1);
  assign Flow_calc_COLUMN_if_and_48_nl = Flow_calc_COLUMN_if_for_10_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[53]);
  assign nl_operator_9_false_acc_102_cse  = conv_u2u_2_3({{1{Flow_calc_COLUMN_if_and_2_psp_54_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_54_sva_1}) + conv_u2u_2_3(signext_2_1(Flow_calc_COLUMN_if_and_48_nl));
  assign Flow_calc_COLUMN_if_and_52_nl = Flow_calc_COLUMN_if_for_8_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[55]);
  assign nl_operator_9_false_acc_62_itm_6_3  = conv_u2u_3_4({{2{Flow_calc_COLUMN_if_and_2_psp_56_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_56_sva_1}) + conv_u2u_3_4(signext_3_1(Flow_calc_COLUMN_if_and_52_nl));
  assign nl_operator_9_false_acc_63_itm_6_3  = conv_u2u_3_4({{2{Flow_calc_COLUMN_if_and_2_psp_58_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_58_sva_1}) + conv_u2u_3_4({{2{Flow_calc_COLUMN_if_and_2_psp_57_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_57_sva_1});
  assign nl_operator_9_false_acc_63_itm_2_1  = conv_u2u_1_2(Flow_calc_COLUMN_if_and_2_psp_58_sva_1)
      + conv_u2u_1_2(Flow_calc_COLUMN_if_and_2_psp_57_sva_1);
  assign Flow_calc_COLUMN_if_and_60_nl = Flow_calc_COLUMN_if_for_4_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[59]);
  assign nl_operator_9_false_acc_64_itm_6_2  = conv_u2u_4_5({{3{Flow_calc_COLUMN_if_and_2_psp_60_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_60_sva_1}) + conv_u2u_4_5(signext_4_1(Flow_calc_COLUMN_if_and_60_nl));
  assign Flow_calc_COLUMN_if_and_1_nl = Flow_calc_COLUMN_if_for_2_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[61]);
  assign nl_operator_9_false_acc_65_itm_6_1  = conv_u2u_5_6({{4{Flow_calc_COLUMN_if_and_seb_1}},
      Flow_calc_COLUMN_if_and_seb_1}) + conv_u2u_5_6(signext_5_1(Flow_calc_COLUMN_if_and_1_nl));
  assign nl_operator_9_false_acc_66_itm_2_0  = conv_u2u_1_3(operator_9_false_asn_76)
      + conv_u2u_2_3({Flow_calc_COLUMN_if_and_2_psp_41_sva_1 , Flow_calc_COLUMN_if_and_2_psp_32_sva_1});
  assign nl_operator_9_false_acc_94_cse  = conv_u2u_1_2(operator_9_false_asn_76)
      + conv_u2u_1_2(Flow_calc_COLUMN_if_and_2_psp_41_sva_1);
  assign nl_operator_9_false_acc_39_itm  = conv_u2u_2_3({Flow_calc_COLUMN_if_and_2_psp_9_sva_1
      , Flow_calc_COLUMN_if_and_2_psp_4_sva_1}) + conv_u2u_2_3({Flow_calc_COLUMN_if_and_2_psp_17_sva_1
      , Flow_calc_COLUMN_if_and_2_psp_8_sva_1});
  assign Flow_calc_COLUMN_if_and_51_nl = Flow_calc_COLUMN_if_for_58_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[5]);
  assign nl_operator_9_false_acc_43_itm_4_1  = conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_39_sva_1
      , ({{1{Flow_calc_COLUMN_if_and_49_seb_1}}, Flow_calc_COLUMN_if_and_49_seb_1})})
      + conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_42_sva_1 , (signext_2_1(Flow_calc_COLUMN_if_and_51_nl))});
  assign nl_operator_9_false_acc_41_itm  = conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_4_sva_1
      , ({{1{Flow_calc_COLUMN_if_and_2_psp_42_sva_1}}, Flow_calc_COLUMN_if_and_2_psp_42_sva_1})})
      + conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_19_sva_1 , ({{1{Flow_calc_COLUMN_if_and_2_psp_34_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_34_sva_1})});
  assign nl_operator_9_false_acc_48_itm  = conv_u2u_5_6({Flow_calc_COLUMN_if_and_2_psp_20_sva_1
      , 1'b0 , Flow_calc_COLUMN_if_and_2_psp_20_sva_1 , 1'b0 , Flow_calc_COLUMN_if_and_2_psp_20_sva_1})
      + conv_u2u_5_6({Flow_calc_COLUMN_if_and_2_psp_21_sva_1 , (signext_4_3({Flow_calc_COLUMN_if_and_2_psp_43_sva_1
      , ({{1{Flow_calc_COLUMN_if_and_2_psp_18_sva_1}}, Flow_calc_COLUMN_if_and_2_psp_18_sva_1})}))});
  assign nl_operator_9_false_acc_44_itm  = conv_u2u_4_5({Flow_calc_COLUMN_if_and_2_psp_9_sva_1
      , ({{2{Flow_calc_COLUMN_if_and_2_psp_38_sva_1}}, Flow_calc_COLUMN_if_and_2_psp_38_sva_1})})
      + conv_u2u_4_5({Flow_calc_COLUMN_if_and_2_psp_10_sva_1 , ({{2{Flow_calc_COLUMN_if_and_2_psp_22_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_22_sva_1})});
  assign Flow_calc_COLUMN_if_and_47_nl = Flow_calc_COLUMN_if_for_56_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[7]);
  assign nl_operator_9_false_acc_45_itm_4_1  = conv_u2u_3_4({Flow_calc_COLUMN_if_and_47_nl
      , ({{1{Flow_calc_COLUMN_if_and_2_psp_37_sva_1}}, Flow_calc_COLUMN_if_and_2_psp_37_sva_1})})
      + conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_8_sva_1 , ({{1{Flow_calc_COLUMN_if_and_2_psp_21_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_21_sva_1})});
  assign Flow_calc_COLUMN_if_and_35_nl = Flow_calc_COLUMN_if_for_50_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[13]);
  assign nl_operator_9_false_acc_52_itm_6_1  = conv_u2u_5_6({Flow_calc_COLUMN_if_and_2_psp_44_sva_1
      , Flow_calc_COLUMN_if_and_2_psp_17_sva_1 , ({{2{Flow_calc_COLUMN_if_and_33_seb_1}},
      Flow_calc_COLUMN_if_and_33_seb_1})}) + conv_u2u_5_6({Flow_calc_COLUMN_if_and_2_psp_45_sva_1
      , Flow_calc_COLUMN_if_and_2_psp_18_sva_1 , (signext_3_1(Flow_calc_COLUMN_if_and_35_nl))});
  assign Flow_calc_COLUMN_if_and_31_nl = Flow_calc_COLUMN_if_for_48_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[15]);
  assign Flow_calc_COLUMN_if_and_39_nl = Flow_calc_COLUMN_if_for_52_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[11]);
  assign nl_operator_9_false_acc_53_itm_6_2  = conv_u2u_4_5({Flow_calc_COLUMN_if_and_2_psp_42_sva_1
      , Flow_calc_COLUMN_if_and_31_nl , ({{1{Flow_calc_COLUMN_if_and_2_psp_12_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_12_sva_1})}) + conv_u2u_4_5({Flow_calc_COLUMN_if_and_2_psp_43_sva_1
      , Flow_calc_COLUMN_if_and_2_psp_16_sva_1 , (signext_2_1(Flow_calc_COLUMN_if_and_39_nl))});
  assign nl_operator_9_false_acc_54_itm_6_3  = conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_38_sva_1
      , ({{1{Flow_calc_COLUMN_if_and_7_seb_1}}, Flow_calc_COLUMN_if_and_7_seb_1})})
      + conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_39_sva_1 , ({{1{Flow_calc_COLUMN_if_and_2_psp_26_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_26_sva_1})});
  assign nl_operator_9_false_acc_55_itm_6_2  = conv_u2u_4_5({Flow_calc_COLUMN_if_and_2_psp_34_sva_1
      , ({{2{Flow_calc_COLUMN_if_and_3_seb_1}}, Flow_calc_COLUMN_if_and_3_seb_1})})
      + conv_u2u_4_5({Flow_calc_COLUMN_if_and_2_psp_35_sva_1 , ({{2{Flow_calc_COLUMN_if_and_2_psp_28_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_28_sva_1})});
  assign Flow_calc_COLUMN_if_and_15_nl = Flow_calc_COLUMN_if_for_40_Flow_calc_COLUMN_if_for_or_1_psp_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[23]);
  assign nl_operator_9_false_acc_56_itm_6_3  = conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_33_sva_1
      , (signext_2_1(Flow_calc_COLUMN_if_and_15_nl))}) + conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_37_sva_1
      , ({{1{Flow_calc_COLUMN_if_and_2_seb_1}}, Flow_calc_COLUMN_if_and_2_seb_1})});
  assign Flow_calc_COLUMN_if_and_4_nl = velocity_value_compare_to_sign_bit_bitwise_OR_complement_35_32_sva_1
      & (Flow_calc_COLUMN_if_acc_6_sdt_sva_1[31]);
  assign nl_operator_9_false_acc_57_itm_6_3  = conv_u2u_3_4({Flow_calc_COLUMN_if_and_4_nl
      , ({{1{Flow_calc_COLUMN_if_and_2_psp_25_sva_1}}, Flow_calc_COLUMN_if_and_2_psp_25_sva_1})})
      + conv_u2u_3_4({Flow_calc_COLUMN_if_and_2_psp_32_sva_1 , ({{1{Flow_calc_COLUMN_if_and_2_psp_24_sva_1}},
      Flow_calc_COLUMN_if_and_2_psp_24_sva_1})});
  assign nl_operator_9_false_acc_109_nl = conv_u2u_3_4(operator_9_false_acc_59_itm_6_4)
      + conv_u2u_3_4(operator_9_false_acc_58_itm_6_4);
  assign operator_9_false_acc_109_nl = nl_operator_9_false_acc_109_nl[3:0];
  assign nl_operator_9_false_acc_110_nl = ({operator_9_false_acc_59_itm_2_1 , Flow_calc_COLUMN_if_and_2_psp_50_sva})
      + conv_u2u_1_3(Flow_calc_COLUMN_if_and_2_psp_48_sva);
  assign operator_9_false_acc_110_nl = nl_operator_9_false_acc_110_nl[2:0];
  assign nl_operator_9_false_acc_84_itm  = conv_u2u_8_9({operator_9_false_acc_109_nl
      , 1'b0 , operator_9_false_acc_110_nl}) + conv_u2u_7_9({operator_9_false_acc_102_cse
      , operator_9_false_acc_102_cse , Flow_calc_COLUMN_if_and_2_psp_54_sva}) + conv_u2u_7_9({operator_9_false_acc_60_itm_6_4
      , operator_9_false_acc_60_itm_3_2 , 1'b0 , Flow_calc_COLUMN_if_and_2_psp_52_sva})
      + conv_u2u_7_9({operator_9_false_acc_65_itm_6_1 , Flow_calc_COLUMN_if_and_seb})
      + conv_u2u_7_9({operator_9_false_acc_64_itm_6_2 , 1'b0 , Flow_calc_COLUMN_if_and_2_psp_60_sva})
      + conv_u2u_7_9({operator_9_false_acc_63_itm_6_3 , operator_9_false_acc_63_itm_2_1
      , Flow_calc_COLUMN_if_and_2_psp_58_sva}) + conv_u2u_7_9({operator_9_false_acc_62_itm_6_3
      , 2'b00 , Flow_calc_COLUMN_if_and_2_psp_56_sva});
  assign nl_operator_9_false_acc_51_nl = conv_u2u_6_7({Flow_calc_COLUMN_if_and_2_psp_46_sva
      , Flow_calc_COLUMN_if_and_2_psp_19_sva , ({{2{Flow_calc_COLUMN_if_and_2_psp_45_sva}},
      Flow_calc_COLUMN_if_and_2_psp_45_sva}) , 1'b1}) + conv_u2u_4_7(operator_9_false_acc_41_itm)
      + conv_u2u_4_7(signext_4_3({Flow_calc_COLUMN_if_and_2_psp_44_sva , ({{1{Flow_calc_COLUMN_if_and_2_psp_10_sva}},
      Flow_calc_COLUMN_if_and_2_psp_10_sva})}));
  assign operator_9_false_acc_51_nl = nl_operator_9_false_acc_51_nl[6:0];
  assign nl_operator_9_false_acc_49_nl = conv_u2s_3_5({Flow_calc_COLUMN_if_and_2_psp_35_sva
      , ({{1{Flow_calc_COLUMN_if_and_57_itm}}, Flow_calc_COLUMN_if_and_57_itm})})
      + conv_s2s_2_5({operator_9_false_acc_40_itm_1 , Flow_calc_COLUMN_if_and_2_psp_16_sva});
  assign operator_9_false_acc_49_nl = nl_operator_9_false_acc_49_nl[4:0];
  assign nl_operator_9_false_acc_69_nl = conv_u2s_5_7({operator_9_false_acc_43_itm_4_1
      , Flow_calc_COLUMN_if_and_49_seb}) + conv_s2s_5_7(operator_9_false_acc_49_nl);
  assign operator_9_false_acc_69_nl = nl_operator_9_false_acc_69_nl[6:0];
  assign nl_operator_9_false_acc_82_nl = conv_u2s_7_9(operator_9_false_acc_51_nl)
      + conv_s2s_7_9(operator_9_false_acc_69_nl);
  assign operator_9_false_acc_82_nl = nl_operator_9_false_acc_82_nl[8:0];
  assign nl_operator_9_false_acc_77_nl = conv_u2u_7_8({operator_9_false_acc_94_cse
      , operator_9_false_acc_94_cse , operator_9_false_acc_66_itm_2_0}) + conv_u2u_6_8({Flow_calc_COLUMN_if_and_2_psp_36_sva
      , 2'b00 , Flow_calc_COLUMN_if_and_2_psp_36_sva , 1'b0 , Flow_calc_COLUMN_if_and_2_psp_36_sva})
      + conv_u2u_5_8({Flow_calc_COLUMN_if_and_2_psp_22_sva , ({{3{Flow_calc_COLUMN_if_and_2_psp_46_sva}},
      Flow_calc_COLUMN_if_and_2_psp_46_sva})}) + conv_u2u_3_8(operator_9_false_acc_39_itm)
      + conv_u2u_3_8({Flow_calc_COLUMN_if_and_55_itm , Flow_calc_COLUMN_if_and_59_itm
      , Flow_calc_COLUMN_if_and_61_itm});
  assign operator_9_false_acc_77_nl = nl_operator_9_false_acc_77_nl[7:0];
  assign nl_operator_9_false_acc_85_itm  = operator_9_false_acc_82_nl + conv_u2s_8_9(operator_9_false_acc_77_nl);
  assign nl_operator_9_false_acc_83_itm  = conv_u2u_7_9({operator_9_false_acc_53_itm_6_2
      , 1'b0 , Flow_calc_COLUMN_if_and_2_psp_12_sva}) + conv_u2u_7_9({operator_9_false_acc_52_itm_6_1
      , Flow_calc_COLUMN_if_and_33_seb}) + conv_u2u_7_9({operator_9_false_acc_57_itm_6_3
      , 1'b0 , Flow_calc_COLUMN_if_and_2_psp_25_sva , Flow_calc_COLUMN_if_and_2_psp_24_sva})
      + conv_u2u_7_9({operator_9_false_acc_56_itm_6_3 , Flow_calc_COLUMN_if_and_2_seb
      , Flow_calc_COLUMN_if_and_2_seb , Flow_calc_COLUMN_if_and_2_seb}) + conv_u2u_7_9({operator_9_false_acc_55_itm_6_2
      , Flow_calc_COLUMN_if_and_3_seb , Flow_calc_COLUMN_if_and_2_psp_28_sva}) +
      conv_u2u_7_9({operator_9_false_acc_54_itm_6_3 , Flow_calc_COLUMN_if_and_7_seb
      , Flow_calc_COLUMN_if_and_2_psp_26_sva , Flow_calc_COLUMN_if_and_2_psp_26_sva})
      + conv_u2u_6_9(operator_9_false_acc_48_itm) + conv_u2u_5_9({operator_9_false_acc_45_itm_4_1
      , Flow_calc_COLUMN_if_and_2_psp_44_sva}) + conv_u2u_5_9(operator_9_false_acc_44_itm);
  assign nl_Flow_calc_COLUMN_acc_itm  = Flow_calc_COLUMN_x_sva + 11'b00000000001;
  assign nl_velocity_value_y_sva  = Flow_calc_COLUMN_if_mul_3_itm - Flow_calc_COLUMN_if_mul_4_itm;
  assign nl_velocity_value_x_sva  = Flow_calc_COLUMN_if_mul_3_itm - Flow_calc_COLUMN_if_mul_2_itm;
  assign nl_Flow_calc_COLUMN_if_if_acc_3_nl = conv_u2s_9_10(Flow_calc_COLUMN_if_if_acc_1_sdt_1[9:1])
      + 10'b1100000001;
  assign Flow_calc_COLUMN_if_if_acc_3_nl = nl_Flow_calc_COLUMN_if_if_acc_3_nl[9:0];
  assign nl_Flow_calc_COLUMN_if_if_acc_nl = conv_s2s_11_12({Flow_calc_COLUMN_if_if_acc_3_nl
      , (Flow_calc_COLUMN_if_if_acc_1_sdt_1[0])}) + conv_s2s_11_12({1'b1 , (~ shift_value_sva)
      , 1'b1});
  assign Flow_calc_COLUMN_if_if_acc_nl = nl_Flow_calc_COLUMN_if_if_acc_nl[11:0];
  assign Flow_calc_COLUMN_if_or_5_nl = (fsm_output[3]) | (fsm_output[6]);
  assign Flow_calc_COLUMN_if_or_6_nl = (fsm_output[5:4]!=2'b00);
  assign Flow_calc_COLUMN_if_mux1h_39_nl = MUX1HOT_v_32_4_2((tensor_shift_value_val_sva_191_96[95:64]),
      (tensor_shift_value_val_sva_191_96[63:32]), (tensor_shift_value_val_sva_191_96[31:0]),
      (tensor_shift_value_val_sva_63_0[31:0]), {Flow_calc_COLUMN_if_or_5_nl , Flow_calc_COLUMN_if_or_6_nl
      , (fsm_output[7]) , (fsm_output[8])});
  assign Flow_calc_COLUMN_if_or_7_nl = (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]);
  assign Flow_calc_COLUMN_if_or_8_nl = (fsm_output[5]) | (fsm_output[8]);
  assign Flow_calc_COLUMN_if_mux1h_40_nl = MUX1HOT_v_32_3_2((tensor_shift_value_val_sva_63_0[31:0]),
      (tensor_shift_value_val_sva_191_96[31:0]), (tensor_shift_value_val_sva_63_0[63:32]),
      {(fsm_output[3]) , Flow_calc_COLUMN_if_or_7_nl , Flow_calc_COLUMN_if_or_8_nl});
  assign nl_mul_sgnd = $signed(Flow_calc_COLUMN_if_mux1h_39_nl) * $signed(Flow_calc_COLUMN_if_mux1h_40_nl);
  assign z_out_1 = $unsigned(nl_mul_sgnd);

  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | (input_1 & {32{sel[1]}});
    result = result | (input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_4_2;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [3:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | (input_1 & {32{sel[1]}});
    result = result | (input_2 & {32{sel[2]}});
    result = result | (input_3 & {32{sel[3]}});
    MUX1HOT_v_32_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | (input_1 & {64{sel[1]}});
    result = result | (input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_13_1_12;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_13_1_12 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input  vector;
  begin
    signext_3_1= {{2{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input  vector;
  begin
    signext_4_1= {{3{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_3;
    input [2:0] vector;
  begin
    signext_4_3= {{1{vector[2]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input  vector;
  begin
    signext_5_1= {{4{vector}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2s_2_5 ;
    input [1:0]  vector ;
  begin
    conv_s2s_2_5 = {{3{vector[1]}}, vector};
  end
  endfunction


  function automatic [6:0] conv_s2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_7 = {{2{vector[4]}}, vector};
  end
  endfunction


  function automatic [8:0] conv_s2s_7_9 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_9 = {{2{vector[6]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_3_5 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_5 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_7 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_7_9 ;
    input [6:0]  vector ;
  begin
    conv_u2s_7_9 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2s_12_13 =  {1'b0, vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_3_8 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_8 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_4_7 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_7 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_5_8 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_8 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_5_9 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_9 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_6_8 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_8 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_6_9 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_9 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_7_9 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_9 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc_struct
// ------------------------------------------------------------------


module OpticalFlow_flow_calc_struct (
  clk, rst, arst_n, tensor_shift_rsc_dat_val, tensor_shift_rsc_vld, tensor_shift_rsc_rdy,
      shift_rsc_dat, shift_rsc_vld, shift_rsc_rdy, output_rsc_dat, output_rsc_vld,
      output_rsc_rdy, widthIn, heightIn, shift_threshold
);
  input clk;
  input rst;
  input arst_n;
  input [191:0] tensor_shift_rsc_dat_val;
  input tensor_shift_rsc_vld;
  output tensor_shift_rsc_rdy;
  input [8:0] shift_rsc_dat;
  input shift_rsc_vld;
  output shift_rsc_rdy;
  output [31:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  input [8:0] shift_threshold;



  // Interconnect Declarations for Component Instantiations 
  OpticalFlow_flow_calc_run OpticalFlow_flow_calc_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_shift_rsc_dat(tensor_shift_rsc_dat_val),
      .tensor_shift_rsc_vld(tensor_shift_rsc_vld),
      .tensor_shift_rsc_rdy(tensor_shift_rsc_rdy),
      .shift_rsc_dat(shift_rsc_dat),
      .shift_rsc_vld(shift_rsc_vld),
      .shift_rsc_rdy(shift_rsc_rdy),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .shift_threshold(shift_threshold)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_flow_calc
// ------------------------------------------------------------------


module OpticalFlow_flow_calc (
  clk, rst, arst_n, tensor_shift_rsc_dat, tensor_shift_rsc_vld, tensor_shift_rsc_rdy,
      shift_rsc_dat, shift_rsc_vld, shift_rsc_rdy, output_rsc_dat, output_rsc_vld,
      output_rsc_rdy, widthIn, heightIn, shift_threshold
);
  input clk;
  input rst;
  input arst_n;
  input [191:0] tensor_shift_rsc_dat;
  input tensor_shift_rsc_vld;
  output tensor_shift_rsc_rdy;
  input [8:0] shift_rsc_dat;
  input shift_rsc_vld;
  output shift_rsc_rdy;
  output [31:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  input [8:0] shift_threshold;



  // Interconnect Declarations for Component Instantiations 
  OpticalFlow_flow_calc_struct OpticalFlow_flow_calc_struct_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_shift_rsc_dat_val(tensor_shift_rsc_dat),
      .tensor_shift_rsc_vld(tensor_shift_rsc_vld),
      .tensor_shift_rsc_rdy(tensor_shift_rsc_rdy),
      .shift_rsc_dat(shift_rsc_dat),
      .shift_rsc_vld(shift_rsc_vld),
      .shift_rsc_rdy(shift_rsc_rdy),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .shift_threshold(shift_threshold)
    );
endmodule




//------> ../OpticalFlow_tensor_weight_x.v4/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Mon Jun 17 23:51:33 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for OpticalFlow_tensor_weight_x_run_run_fsm_1
  parameter
    main_C_0 = 1'd0,
    main_C_1 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : OpticalFlow_tensor_weight_x_run_run_fsm_1
    case (state_var)
      main_C_1 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_1;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_staller
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_staller (
  run_wen, tensor_y_rsci_wen_comp, tensor_shift_rsci_wen_comp, shift_rsci_wen_comp
);
  output run_wen;
  input tensor_y_rsci_wen_comp;
  input tensor_shift_rsci_wen_comp;
  input shift_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = tensor_y_rsci_wen_comp & tensor_shift_rsci_wen_comp & shift_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_wait_dp (
  clk, rst, arst_n, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z,
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z, Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z,
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z, run_wen, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg, Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg,
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg, Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg
);
  input clk;
  input rst;
  input arst_n;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z;
  input [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z;
  input [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z;
  input [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z;
  input run_wen;
  output [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg;
  output [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg;
  output [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg;
  output [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg;
  output [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg;
  output [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg;
  output [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg;
  reg [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg;
  output [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg;
  reg [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg;
  output [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg;
  reg [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg;



  // Interconnect Declarations for Component Instantiations 
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg <= Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg <= Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg <= Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg <= Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg <= Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg <= Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg <= Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg <= Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg <= Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_shift_rsci_shift_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_shift_rsci_shift_wait_dp (
  clk, rst, arst_n, shift_rsci_oswt, shift_rsci_wen_comp, shift_rsci_biwt, shift_rsci_bdwt,
      shift_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input shift_rsci_oswt;
  output shift_rsci_wen_comp;
  input shift_rsci_biwt;
  input shift_rsci_bdwt;
  output shift_rsci_bcwt;
  reg shift_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign shift_rsci_wen_comp = (~ shift_rsci_oswt) | shift_rsci_biwt | shift_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      shift_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      shift_rsci_bcwt <= 1'b0;
    end
    else begin
      shift_rsci_bcwt <= ~((~(shift_rsci_bcwt | shift_rsci_biwt)) | shift_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_shift_rsci_shift_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_shift_rsci_shift_wait_ctrl (
  run_wen, shift_rsci_oswt, shift_rsci_biwt, shift_rsci_bdwt, shift_rsci_bcwt, shift_rsci_irdy,
      shift_rsci_ivld_run_sct
);
  input run_wen;
  input shift_rsci_oswt;
  output shift_rsci_biwt;
  output shift_rsci_bdwt;
  input shift_rsci_bcwt;
  input shift_rsci_irdy;
  output shift_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire shift_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign shift_rsci_bdwt = shift_rsci_oswt & run_wen;
  assign shift_rsci_biwt = shift_rsci_ogwt & shift_rsci_irdy;
  assign shift_rsci_ogwt = shift_rsci_oswt & (~ shift_rsci_bcwt);
  assign shift_rsci_ivld_run_sct = shift_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_tensor_shift_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_tensor_shift_wait_dp (
  clk, rst, arst_n, tensor_shift_rsci_oswt, tensor_shift_rsci_wen_comp, tensor_shift_rsci_biwt,
      tensor_shift_rsci_bdwt, tensor_shift_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input tensor_shift_rsci_oswt;
  output tensor_shift_rsci_wen_comp;
  input tensor_shift_rsci_biwt;
  input tensor_shift_rsci_bdwt;
  output tensor_shift_rsci_bcwt;
  reg tensor_shift_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign tensor_shift_rsci_wen_comp = (~ tensor_shift_rsci_oswt) | tensor_shift_rsci_biwt
      | tensor_shift_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      tensor_shift_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      tensor_shift_rsci_bcwt <= 1'b0;
    end
    else begin
      tensor_shift_rsci_bcwt <= ~((~(tensor_shift_rsci_bcwt | tensor_shift_rsci_biwt))
          | tensor_shift_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_tensor_shift_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_tensor_shift_wait_ctrl (
  run_wen, tensor_shift_rsci_oswt, tensor_shift_rsci_biwt, tensor_shift_rsci_bdwt,
      tensor_shift_rsci_bcwt, tensor_shift_rsci_irdy, tensor_shift_rsci_ivld_run_sct
);
  input run_wen;
  input tensor_shift_rsci_oswt;
  output tensor_shift_rsci_biwt;
  output tensor_shift_rsci_bdwt;
  input tensor_shift_rsci_bcwt;
  input tensor_shift_rsci_irdy;
  output tensor_shift_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire tensor_shift_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign tensor_shift_rsci_bdwt = tensor_shift_rsci_oswt & run_wen;
  assign tensor_shift_rsci_biwt = tensor_shift_rsci_ogwt & tensor_shift_rsci_irdy;
  assign tensor_shift_rsci_ogwt = tensor_shift_rsci_oswt & (~ tensor_shift_rsci_bcwt);
  assign tensor_shift_rsci_ivld_run_sct = tensor_shift_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_tensor_y_rsci_tensor_y_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_tensor_y_rsci_tensor_y_wait_ctrl (
  run_wen, tensor_y_rsci_iswt0, tensor_y_rsci_irdy_run_sct
);
  input run_wen;
  input tensor_y_rsci_iswt0;
  output tensor_y_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign tensor_y_rsci_irdy_run_sct = tensor_y_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_shift_rsci
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_shift_rsci (
  clk, rst, arst_n, shift_rsc_dat, shift_rsc_vld, shift_rsc_rdy, run_wen, shift_rsci_oswt,
      shift_rsci_wen_comp, shift_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [8:0] shift_rsc_dat;
  output shift_rsc_vld;
  input shift_rsc_rdy;
  input run_wen;
  input shift_rsci_oswt;
  output shift_rsci_wen_comp;
  input [8:0] shift_rsci_idat;


  // Interconnect Declarations
  wire shift_rsci_biwt;
  wire shift_rsci_bdwt;
  wire shift_rsci_bcwt;
  wire shift_rsci_irdy;
  wire shift_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd9)) shift_rsci (
      .irdy(shift_rsci_irdy),
      .ivld(shift_rsci_ivld_run_sct),
      .idat(shift_rsci_idat),
      .rdy(shift_rsc_rdy),
      .vld(shift_rsc_vld),
      .dat(shift_rsc_dat)
    );
  OpticalFlow_tensor_weight_x_run_shift_rsci_shift_wait_ctrl OpticalFlow_tensor_weight_x_run_shift_rsci_shift_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .shift_rsci_oswt(shift_rsci_oswt),
      .shift_rsci_biwt(shift_rsci_biwt),
      .shift_rsci_bdwt(shift_rsci_bdwt),
      .shift_rsci_bcwt(shift_rsci_bcwt),
      .shift_rsci_irdy(shift_rsci_irdy),
      .shift_rsci_ivld_run_sct(shift_rsci_ivld_run_sct)
    );
  OpticalFlow_tensor_weight_x_run_shift_rsci_shift_wait_dp OpticalFlow_tensor_weight_x_run_shift_rsci_shift_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .shift_rsci_oswt(shift_rsci_oswt),
      .shift_rsci_wen_comp(shift_rsci_wen_comp),
      .shift_rsci_biwt(shift_rsci_biwt),
      .shift_rsci_bdwt(shift_rsci_bdwt),
      .shift_rsci_bcwt(shift_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_tensor_shift_rsci
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_tensor_shift_rsci (
  clk, rst, arst_n, tensor_shift_rsc_dat, tensor_shift_rsc_vld, tensor_shift_rsc_rdy,
      run_wen, tensor_shift_rsci_oswt, tensor_shift_rsci_wen_comp, tensor_shift_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [191:0] tensor_shift_rsc_dat;
  output tensor_shift_rsc_vld;
  input tensor_shift_rsc_rdy;
  input run_wen;
  input tensor_shift_rsci_oswt;
  output tensor_shift_rsci_wen_comp;
  input [191:0] tensor_shift_rsci_idat;


  // Interconnect Declarations
  wire tensor_shift_rsci_biwt;
  wire tensor_shift_rsci_bdwt;
  wire tensor_shift_rsci_bcwt;
  wire tensor_shift_rsci_irdy;
  wire tensor_shift_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd192)) tensor_shift_rsci (
      .irdy(tensor_shift_rsci_irdy),
      .ivld(tensor_shift_rsci_ivld_run_sct),
      .idat(tensor_shift_rsci_idat),
      .rdy(tensor_shift_rsc_rdy),
      .vld(tensor_shift_rsc_vld),
      .dat(tensor_shift_rsc_dat)
    );
  OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_tensor_shift_wait_ctrl OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_tensor_shift_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .tensor_shift_rsci_oswt(tensor_shift_rsci_oswt),
      .tensor_shift_rsci_biwt(tensor_shift_rsci_biwt),
      .tensor_shift_rsci_bdwt(tensor_shift_rsci_bdwt),
      .tensor_shift_rsci_bcwt(tensor_shift_rsci_bcwt),
      .tensor_shift_rsci_irdy(tensor_shift_rsci_irdy),
      .tensor_shift_rsci_ivld_run_sct(tensor_shift_rsci_ivld_run_sct)
    );
  OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_tensor_shift_wait_dp OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_tensor_shift_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_shift_rsci_oswt(tensor_shift_rsci_oswt),
      .tensor_shift_rsci_wen_comp(tensor_shift_rsci_wen_comp),
      .tensor_shift_rsci_biwt(tensor_shift_rsci_biwt),
      .tensor_shift_rsci_bdwt(tensor_shift_rsci_bdwt),
      .tensor_shift_rsci_bcwt(tensor_shift_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run_tensor_y_rsci
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run_tensor_y_rsci (
  tensor_y_rsc_dat, tensor_y_rsc_vld, tensor_y_rsc_rdy, run_wen, tensor_y_rsci_oswt,
      tensor_y_rsci_wen_comp, tensor_y_rsci_idat_mxwt
);
  input [383:0] tensor_y_rsc_dat;
  input tensor_y_rsc_vld;
  output tensor_y_rsc_rdy;
  input run_wen;
  input tensor_y_rsci_oswt;
  output tensor_y_rsci_wen_comp;
  output [383:0] tensor_y_rsci_idat_mxwt;


  // Interconnect Declarations
  wire tensor_y_rsci_irdy_run_sct;
  wire tensor_y_rsci_ivld;
  wire [383:0] tensor_y_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd1),
  .width(32'sd384)) tensor_y_rsci (
      .rdy(tensor_y_rsc_rdy),
      .vld(tensor_y_rsc_vld),
      .dat(tensor_y_rsc_dat),
      .irdy(tensor_y_rsci_irdy_run_sct),
      .ivld(tensor_y_rsci_ivld),
      .idat(tensor_y_rsci_idat)
    );
  OpticalFlow_tensor_weight_x_run_tensor_y_rsci_tensor_y_wait_ctrl OpticalFlow_tensor_weight_x_run_tensor_y_rsci_tensor_y_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .tensor_y_rsci_iswt0(tensor_y_rsci_oswt),
      .tensor_y_rsci_irdy_run_sct(tensor_y_rsci_irdy_run_sct)
    );
  assign tensor_y_rsci_idat_mxwt = tensor_y_rsci_idat;
  assign tensor_y_rsci_wen_comp = (~ tensor_y_rsci_oswt) | tensor_y_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_run
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_run (
  clk, rst, arst_n, tensor_y_rsc_dat, tensor_y_rsc_vld, tensor_y_rsc_rdy, tensor_shift_rsc_dat,
      tensor_shift_rsc_vld, tensor_shift_rsc_rdy, shift_rsc_dat, shift_rsc_vld, shift_rsc_rdy,
      widthIn, heightIn, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z,
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b, Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z,
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b, Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z,
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b, Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z,
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b, Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z
);
  input clk;
  input rst;
  input arst_n;
  input [383:0] tensor_y_rsc_dat;
  input tensor_y_rsc_vld;
  output tensor_y_rsc_rdy;
  output [191:0] tensor_shift_rsc_dat;
  output tensor_shift_rsc_vld;
  input tensor_shift_rsc_rdy;
  output [8:0] shift_rsc_dat;
  output shift_rsc_vld;
  input shift_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  output [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b;
  reg [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z;
  output [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b;
  reg [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z;
  output [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b;
  reg [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z;
  output [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b;
  reg [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z;
  output [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b;
  reg [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z;
  output [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b;
  reg [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b;
  input [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z;
  output [63:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b;
  reg [63:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b;
  input [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z;
  output [63:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b;
  reg [63:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b;
  input [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z;
  output [63:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b;
  reg [63:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b;
  input [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z;


  // Interconnect Declarations
  wire run_wen;
  wire tensor_y_rsci_wen_comp;
  wire [383:0] tensor_y_rsci_idat_mxwt;
  wire tensor_shift_rsci_wen_comp;
  wire shift_rsci_wen_comp;
  reg [8:0] shift_rsci_idat;
  wire [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg;
  wire [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg;
  wire [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg;
  wire [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg;
  wire [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg;
  wire [93:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg;
  wire [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg;
  wire [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg;
  wire [92:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg;
  reg [31:0] tensor_shift_rsci_idat_191_160;
  reg [31:0] tensor_shift_rsci_idat_159_128;
  reg [31:0] tensor_shift_rsci_idat_127_96;
  reg [31:0] tensor_shift_rsci_idat_95_64;
  reg [31:0] tensor_shift_rsci_idat_63_32;
  reg [31:0] tensor_shift_rsci_idat_31_0;
  wire [1:0] fsm_output;
  wire [9:0] operator_9_false_1_acc_tmp;
  wire [10:0] nl_operator_9_false_1_acc_tmp;
  wire Tensor_weight_x_COLUMN_equal_tmp;
  wire or_tmp_3;
  wire or_tmp_35;
  wire or_tmp_36;
  reg operator_9_false_acc_76_itm_1_0;
  reg main_stage_0_2;
  reg Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_3;
  reg main_stage_0_4;
  reg Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_2;
  reg main_stage_0_3;
  reg Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_1;
  reg operator_11_false_1_slc_operator_11_false_1_acc_11_itm_3;
  reg exitL_exit_Tensor_weight_x_ROW_sva;
  reg Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_4;
  reg [10:0] Tensor_weight_x_COLUMN_x_lpi_1_dfm;
  wire exit_Tensor_weight_x_ROW_sva_2_mx0w0;
  reg reg_shift_rsci_oswt_cse;
  wire Tensor_weight_x_COLUMN_if_1_and_95_cse;
  wire tensor0_val_and_cse;
  reg reg_tensor_y_rsci_oswt_cse;
  wire tensor_buf0_val_and_cse;
  wire and_184_cse;
  wire [95:0] Tensor_weight_x_COLUMN_if_1_lshift_3_itm;
  wire [95:0] z_out;
  wire [95:0] z_out_1;
  wire [8:0] z_out_2;
  wire [9:0] nl_z_out_2;
  reg [63:0] tensor_buf1_val_255_192_lpi_1;
  reg [63:0] tensor_buf1_val_127_64_lpi_1;
  reg [63:0] tensor_buf1_val_63_0_lpi_1;
  reg [8:0] Tensor_weight_x_ROW_y_lpi_1_dfm;
  reg [63:0] tensor_buf0_val_383_320_lpi_1_dfm;
  reg [63:0] tensor_buf0_val_191_128_lpi_1_dfm;
  reg [63:0] tensor_buf0_val_127_64_lpi_1_dfm;
  reg [94:0] Tensor_weight_x_COLUMN_if_1_acc_psp_sva;
  reg [94:0] Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_64_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_63_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_62_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_61_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_60_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_59_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_58_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_57_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_56_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_55_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_54_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_53_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_52_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_51_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_50_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_49_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_48_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_47_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_46_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_45_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_44_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_43_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_42_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_41_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_40_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_39_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_38_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_37_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_36_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_35_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_34_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_33_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_32_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_31_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_30_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_29_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_28_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_27_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_26_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_25_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_24_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_23_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_22_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_21_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_20_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_19_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_18_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_17_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_16_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_15_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_14_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_13_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_12_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_9_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_8_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_7_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_6_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_5_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_4_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_3_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_2_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_1_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_80_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_79_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_78_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_77_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_76_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_75_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_74_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_73_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_72_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_71_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_70_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_69_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_68_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_67_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_66_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_65_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_88_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_87_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_86_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_85_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_84_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_83_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_82_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_81_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_92_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_91_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_90_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_89_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_94_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_93_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg Tensor_weight_x_COLUMN_if_1_for_95_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva;
  reg [31:0] Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm;
  reg [63:0] tensor0_val_0_lpi_1_dfm_1;
  reg [63:0] tensor0_val_1_lpi_1_dfm_1;
  reg [63:0] tensor0_val_2_lpi_1_dfm_1;
  reg [63:0] tensor0_val_3_lpi_1_dfm_1;
  reg [63:0] tensor0_val_4_lpi_1_dfm_1;
  reg [94:0] Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1;
  reg [94:0] Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1;
  reg [8:0] Tensor_weight_x_COLUMN_if_1_ac_int_cctor_1_sva_1;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_asn_28_itm_1;
  reg [8:0] operator_9_false_acc_105_itm_1;
  wire [10:0] nl_operator_9_false_acc_105_itm_1;
  reg [8:0] operator_9_false_acc_104_itm_1;
  wire [9:0] nl_operator_9_false_acc_104_itm_1;
  reg [8:0] operator_9_false_acc_103_itm_1;
  reg [8:0] operator_9_false_acc_102_itm_1;
  reg [5:0] operator_9_false_acc_79_itm_1;
  wire [6:0] nl_operator_9_false_acc_79_itm_1;
  reg [5:0] operator_9_false_acc_68_itm_1;
  wire [6:0] nl_operator_9_false_acc_68_itm_1;
  reg [5:0] operator_9_false_acc_71_itm_1;
  wire [7:0] nl_operator_9_false_acc_71_itm_1;
  reg [5:0] operator_9_false_acc_70_itm_1;
  wire [7:0] nl_operator_9_false_acc_70_itm_1;
  reg [6:0] operator_9_false_acc_78_itm_1;
  wire [8:0] nl_operator_9_false_acc_78_itm_1;
  reg [6:0] operator_9_false_acc_77_itm_1;
  wire [8:0] nl_operator_9_false_acc_77_itm_1;
  reg [6:0] operator_9_false_acc_75_itm_1;
  wire [8:0] nl_operator_9_false_acc_75_itm_1;
  reg [7:0] operator_9_false_acc_97_itm_1;
  wire [9:0] nl_operator_9_false_acc_97_itm_1;
  reg [8:0] operator_9_false_acc_108_itm_1;
  wire [9:0] nl_operator_9_false_acc_108_itm_1;
  reg [8:0] operator_9_false_acc_107_itm_1;
  wire [9:0] nl_operator_9_false_acc_107_itm_1;
  reg [31:0] Tensor_weight_x_COLUMN_if_1_slc_95_64_5_itm_1;
  reg [31:0] Tensor_weight_x_COLUMN_if_1_slc_95_64_4_itm_1;
  reg [31:0] Tensor_weight_x_COLUMN_if_1_slc_95_64_3_itm_1;
  reg [63:0] Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_10_itm_1;
  reg [31:0] Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm_1;
  reg operator_11_false_1_slc_operator_11_false_1_acc_11_itm_1;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_94_1;
  wire [94:0] nl_Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_94_1;
  reg Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_0;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_94_1;
  wire [94:0] nl_Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_94_1;
  reg Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_0;
  reg Tensor_weight_x_COLUMN_if_1_acc_16_itm_1_0;
  reg [6:0] operator_9_false_acc_81_itm_1_7_1;
  wire [7:0] nl_operator_9_false_acc_81_itm_1_7_1;
  reg [5:0] operator_9_false_acc_76_itm_1_6_1;
  wire [7:0] nl_operator_9_false_acc_76_itm_1_6_1;
  reg [1:0] operator_9_false_acc_74_itm_1_6_5;
  wire [2:0] nl_operator_9_false_acc_74_itm_1_6_5;
  reg [2:0] operator_9_false_acc_74_itm_1_2_0;
  wire [3:0] nl_operator_9_false_acc_74_itm_1_2_0;
  reg [1:0] operator_9_false_acc_96_itm_1_7_6;
  wire [2:0] nl_operator_9_false_acc_96_itm_1_7_6;
  reg [4:0] operator_9_false_acc_106_itm_1_8_4;
  wire [6:0] nl_operator_9_false_acc_106_itm_1_8_4;
  reg [3:0] operator_9_false_acc_106_itm_1_3_0;
  wire [4:0] nl_operator_9_false_acc_106_itm_1_3_0;
  wire exitL_exit_Tensor_weight_x_ROW_sva_mx0;
  wire [10:0] Tensor_weight_x_COLUMN_x_lpi_1_dfm_mx0w0;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_34_sva_1;
  wire [94:0] Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1;
  wire [95:0] nl_Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1;
  wire [94:0] Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1;
  wire [95:0] nl_Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1;
  wire [94:0] Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1;
  wire [95:0] nl_Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1;
  wire [94:0] Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1;
  wire [96:0] nl_Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1;
  wire [94:0] Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1;
  wire [96:0] nl_Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_68_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_72_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_70_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_51_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_66_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_50_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_67_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_49_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_69_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_48_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_83_sva_1;
  wire [94:0] Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1;
  wire [95:0] nl_Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_54_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_82_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_64_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_53_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_65_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_52_sva_1;
  wire [1:0] operator_9_false_acc_138_cse_1;
  wire [2:0] nl_operator_9_false_acc_138_cse_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_84_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_73_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_81_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_32_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_44_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_43_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_psp_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_24_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_45_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_46_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_28_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_41_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_8_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_86_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_76_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_18_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_19_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_35_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_90_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_36_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_22_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_79_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_77_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_85_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_75_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_17_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_12_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_21_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_65_seb_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_87_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_88_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_42_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_78_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_16_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_10_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_39_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_71_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_74_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_9_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_38_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_20_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_37_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_92_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_33_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_4_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_89_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_1_psp_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_26_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_25_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_91_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_57_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_56_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_60_sva_1;
  wire Tensor_weight_x_COLUMN_if_1_and_34_seb_1;
  wire Tensor_weight_x_COLUMN_if_1_and_2_psp_58_sva_1;
  wire operator_9_false_asn_221;
  reg Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_94;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_93_0;
  reg Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_94;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_93_0;
  reg Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_94;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_93_0;
  wire [8:0] Tensor_weight_x_COLUMN_if_1_mux_17_cse;
  reg Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_94;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_93_0;
  reg Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_94;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_93_0;
  reg Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_94;
  reg [93:0] Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_93_0;
  wire Tensor_weight_x_COLUMN_if_1_and_105_cse;
  wire operator_11_false_acc_itm_11_1;

  wire Tensor_weight_x_COLUMN_if_1_not_9_nl;
  wire Tensor_weight_x_COLUMN_if_1_not_10_nl;
  wire Tensor_weight_x_COLUMN_if_1_not_11_nl;
  wire Tensor_weight_x_COLUMN_if_1_not_12_nl;
  wire Tensor_weight_x_COLUMN_if_1_not_13_nl;
  wire Tensor_weight_x_COLUMN_if_1_not_14_nl;
  wire Tensor_weight_x_COLUMN_if_1_not_15_nl;
  wire[63:0] Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_9_nl;
  wire Tensor_weight_x_ROW_not_46_nl;
  wire[63:0] Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_11_nl;
  wire Tensor_weight_x_ROW_not_47_nl;
  wire[63:0] Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_8_nl;
  wire Tensor_weight_x_ROW_not_45_nl;
  wire[63:0] Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_7_nl;
  wire Tensor_weight_x_ROW_not_44_nl;
  wire[63:0] Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_12_nl;
  wire Tensor_weight_x_ROW_not_48_nl;
  wire[63:0] or_nl;
  wire nor_1_nl;
  wire nor_nl;
  wire[63:0] Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_2_nl;
  wire Tensor_weight_x_ROW_not_38_nl;
  wire[63:0] Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_3_nl;
  wire Tensor_weight_x_ROW_not_41_nl;
  wire[11:0] Tensor_weight_x_COLUMN_aelse_acc_nl;
  wire[12:0] nl_Tensor_weight_x_COLUMN_aelse_acc_nl;
  wire Tensor_weight_x_ROW_not_42_nl;
  wire[63:0] Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_5_nl;
  wire Tensor_weight_x_ROW_not_40_nl;
  wire[3:0] operator_9_false_acc_135_nl;
  wire[4:0] nl_operator_9_false_acc_135_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_47_nl;
  wire[1:0] operator_9_false_acc_141_nl;
  wire[2:0] nl_operator_9_false_acc_141_nl;
  wire[2:0] operator_9_false_acc_142_nl;
  wire[3:0] nl_operator_9_false_acc_142_nl;
  wire[3:0] operator_9_false_acc_143_nl;
  wire[4:0] nl_operator_9_false_acc_143_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_36_nl;
  wire[3:0] operator_9_false_acc_144_nl;
  wire[4:0] nl_operator_9_false_acc_144_nl;
  wire[3:0] operator_9_false_acc_145_nl;
  wire[4:0] nl_operator_9_false_acc_145_nl;
  wire[1:0] operator_9_false_acc_146_nl;
  wire[2:0] nl_operator_9_false_acc_146_nl;
  wire[3:0] operator_9_false_acc_120_nl;
  wire[4:0] nl_operator_9_false_acc_120_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_4_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_32_nl;
  wire[4:0] operator_9_false_acc_121_nl;
  wire[5:0] nl_operator_9_false_acc_121_nl;
  wire[4:0] operator_9_false_acc_122_nl;
  wire[5:0] nl_operator_9_false_acc_122_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_20_nl;
  wire[8:0] operator_9_false_acc_nl;
  wire[9:0] nl_operator_9_false_acc_nl;
  wire[8:0] operator_9_false_acc_117_nl;
  wire[10:0] nl_operator_9_false_acc_117_nl;
  wire[8:0] operator_9_false_acc_119_nl;
  wire[9:0] nl_operator_9_false_acc_119_nl;
  wire[8:0] operator_9_false_acc_116_nl;
  wire[9:0] nl_operator_9_false_acc_116_nl;
  wire[8:0] operator_9_false_acc_111_nl;
  wire[9:0] nl_operator_9_false_acc_111_nl;
  wire[7:0] operator_9_false_acc_101_nl;
  wire[8:0] nl_operator_9_false_acc_101_nl;
  wire[7:0] operator_9_false_acc_100_nl;
  wire[9:0] nl_operator_9_false_acc_100_nl;
  wire[8:0] operator_9_false_acc_110_nl;
  wire[10:0] nl_operator_9_false_acc_110_nl;
  wire[8:0] operator_9_false_acc_103_nl;
  wire[10:0] nl_operator_9_false_acc_103_nl;
  wire[5:0] operator_9_false_acc_123_nl;
  wire[6:0] nl_operator_9_false_acc_123_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_28_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_31_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_39_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_33_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_35_nl;
  wire[8:0] operator_9_false_acc_118_nl;
  wire[11:0] nl_operator_9_false_acc_118_nl;
  wire[8:0] operator_9_false_acc_102_nl;
  wire[10:0] nl_operator_9_false_acc_102_nl;
  wire[4:0] operator_9_false_acc_124_nl;
  wire[5:0] nl_operator_9_false_acc_124_nl;
  wire[1:0] operator_9_false_acc_125_nl;
  wire[2:0] nl_operator_9_false_acc_125_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_89_nl;
  wire[4:0] operator_9_false_acc_56_nl;
  wire[6:0] nl_operator_9_false_acc_56_nl;
  wire[4:0] operator_9_false_acc_69_nl;
  wire[5:0] nl_operator_9_false_acc_69_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_79_nl;
  wire[3:0] operator_9_false_acc_127_nl;
  wire[4:0] nl_operator_9_false_acc_127_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_83_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_81_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_87_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_63_nl;
  wire[3:0] operator_9_false_acc_128_nl;
  wire[4:0] nl_operator_9_false_acc_128_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_71_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_67_nl;
  wire[10:0] operator_11_false_acc_nl;
  wire[11:0] nl_operator_11_false_acc_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_91_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_93_nl;
  wire Tensor_weight_x_ROW_not_43_nl;
  wire[8:0] Tensor_weight_x_COLUMN_if_2_mux_nl;
  wire[8:0] Tensor_weight_x_ROW_acc_nl;
  wire[9:0] nl_Tensor_weight_x_ROW_acc_nl;
  wire Tensor_weight_x_ROW_not_34_nl;
  wire[94:0] Tensor_weight_x_COLUMN_if_1_acc_4_nl;
  wire[96:0] nl_Tensor_weight_x_COLUMN_if_1_acc_4_nl;
  wire[93:0] Tensor_weight_x_COLUMN_if_1_acc_22_nl;
  wire[94:0] nl_Tensor_weight_x_COLUMN_if_1_acc_22_nl;
  wire Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_nl;
  wire Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_nl;
  wire[11:0] operator_11_false_1_acc_nl;
  wire[12:0] nl_operator_11_false_1_acc_nl;
  wire[11:0] operator_11_false_acc_nl_1;
  wire[12:0] nl_operator_11_false_acc_nl_1;
  wire[10:0] Tensor_weight_x_COLUMN_if_2_mux_1_nl;
  wire[10:0] Tensor_weight_x_COLUMN_acc_1_nl;
  wire[11:0] nl_Tensor_weight_x_COLUMN_acc_1_nl;
  wire Tensor_weight_x_ROW_Tensor_weight_x_ROW_Tensor_weight_x_ROW_Tensor_weight_x_ROW_not_nl;
  wire Tensor_weight_x_COLUMN_if_1_and_70_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [95:0] nl_Tensor_weight_x_COLUMN_if_1_lshift_3_rg_a;
  assign nl_Tensor_weight_x_COLUMN_if_1_lshift_3_rg_a = {Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_94
      , Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_93_0 , 1'b0};
  wire Tensor_weight_x_COLUMN_if_1_mux_20_nl;
  wire[93:0] Tensor_weight_x_COLUMN_if_1_mux_23_nl;
  wire [95:0] nl_Tensor_weight_x_COLUMN_if_1_lshift_rg_a;
  assign Tensor_weight_x_COLUMN_if_1_mux_20_nl = MUX_s_1_2_2((Tensor_weight_x_COLUMN_if_1_acc_psp_sva[94]),
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_94, fsm_output[1]);
  assign Tensor_weight_x_COLUMN_if_1_mux_23_nl = MUX_v_94_2_2((Tensor_weight_x_COLUMN_if_1_acc_psp_sva[93:0]),
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_93_0, fsm_output[1]);
  assign nl_Tensor_weight_x_COLUMN_if_1_lshift_rg_a = {Tensor_weight_x_COLUMN_if_1_mux_20_nl
      , Tensor_weight_x_COLUMN_if_1_mux_23_nl , 1'b0};
  wire Tensor_weight_x_COLUMN_if_1_mux_18_nl;
  wire[93:0] Tensor_weight_x_COLUMN_if_1_mux_24_nl;
  wire [95:0] nl_Tensor_weight_x_COLUMN_if_1_lshift_1_rg_a;
  assign Tensor_weight_x_COLUMN_if_1_mux_18_nl = MUX_s_1_2_2((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva[94]),
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_94, fsm_output[1]);
  assign Tensor_weight_x_COLUMN_if_1_mux_24_nl = MUX_v_94_2_2((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva[93:0]),
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_93_0, fsm_output[1]);
  assign nl_Tensor_weight_x_COLUMN_if_1_lshift_1_rg_a = {Tensor_weight_x_COLUMN_if_1_mux_18_nl
      , Tensor_weight_x_COLUMN_if_1_mux_24_nl , 1'b0};
  wire [191:0] nl_OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_inst_tensor_shift_rsci_idat;
  assign nl_OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_inst_tensor_shift_rsci_idat
      = {tensor_shift_rsci_idat_191_160 , tensor_shift_rsci_idat_159_128 , tensor_shift_rsci_idat_127_96
      , tensor_shift_rsci_idat_95_64 , tensor_shift_rsci_idat_63_32 , tensor_shift_rsci_idat_31_0};
  mgc_shift_l_v5 #(.width_a(32'sd96),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd96)) Tensor_weight_x_COLUMN_if_1_lshift_3_rg (
      .a(nl_Tensor_weight_x_COLUMN_if_1_lshift_3_rg_a[95:0]),
      .s(z_out_2),
      .z(Tensor_weight_x_COLUMN_if_1_lshift_3_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd96),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd96)) Tensor_weight_x_COLUMN_if_1_lshift_rg (
      .a(nl_Tensor_weight_x_COLUMN_if_1_lshift_rg_a[95:0]),
      .s(Tensor_weight_x_COLUMN_if_1_mux_17_cse),
      .z(z_out)
    );
  mgc_shift_l_v5 #(.width_a(32'sd96),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd96)) Tensor_weight_x_COLUMN_if_1_lshift_1_rg (
      .a(nl_Tensor_weight_x_COLUMN_if_1_lshift_1_rg_a[95:0]),
      .s(Tensor_weight_x_COLUMN_if_1_mux_17_cse),
      .z(z_out_1)
    );
  OpticalFlow_tensor_weight_x_run_tensor_y_rsci OpticalFlow_tensor_weight_x_run_tensor_y_rsci_inst
      (
      .tensor_y_rsc_dat(tensor_y_rsc_dat),
      .tensor_y_rsc_vld(tensor_y_rsc_vld),
      .tensor_y_rsc_rdy(tensor_y_rsc_rdy),
      .run_wen(run_wen),
      .tensor_y_rsci_oswt(reg_tensor_y_rsci_oswt_cse),
      .tensor_y_rsci_wen_comp(tensor_y_rsci_wen_comp),
      .tensor_y_rsci_idat_mxwt(tensor_y_rsci_idat_mxwt)
    );
  OpticalFlow_tensor_weight_x_run_tensor_shift_rsci OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_shift_rsc_dat(tensor_shift_rsc_dat),
      .tensor_shift_rsc_vld(tensor_shift_rsc_vld),
      .tensor_shift_rsc_rdy(tensor_shift_rsc_rdy),
      .run_wen(run_wen),
      .tensor_shift_rsci_oswt(reg_shift_rsci_oswt_cse),
      .tensor_shift_rsci_wen_comp(tensor_shift_rsci_wen_comp),
      .tensor_shift_rsci_idat(nl_OpticalFlow_tensor_weight_x_run_tensor_shift_rsci_inst_tensor_shift_rsci_idat[191:0])
    );
  OpticalFlow_tensor_weight_x_run_shift_rsci OpticalFlow_tensor_weight_x_run_shift_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .shift_rsc_dat(shift_rsc_dat),
      .shift_rsc_vld(shift_rsc_vld),
      .shift_rsc_rdy(shift_rsc_rdy),
      .run_wen(run_wen),
      .shift_rsci_oswt(reg_shift_rsci_oswt_cse),
      .shift_rsci_wen_comp(shift_rsci_wen_comp),
      .shift_rsci_idat(shift_rsci_idat)
    );
  OpticalFlow_tensor_weight_x_run_wait_dp OpticalFlow_tensor_weight_x_run_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z),
      .run_wen(run_wen),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg)
    );
  OpticalFlow_tensor_weight_x_run_staller OpticalFlow_tensor_weight_x_run_staller_inst
      (
      .run_wen(run_wen),
      .tensor_y_rsci_wen_comp(tensor_y_rsci_wen_comp),
      .tensor_shift_rsci_wen_comp(tensor_shift_rsci_wen_comp),
      .shift_rsci_wen_comp(shift_rsci_wen_comp)
    );
  OpticalFlow_tensor_weight_x_run_run_fsm OpticalFlow_tensor_weight_x_run_run_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign Tensor_weight_x_COLUMN_if_1_and_95_cse = run_wen & ((Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_4
      & exitL_exit_Tensor_weight_x_ROW_sva & (fsm_output[0])) | or_tmp_3);
  assign Tensor_weight_x_COLUMN_if_1_and_105_cse = run_wen & (fsm_output[1]);
  assign tensor0_val_and_cse = run_wen & ((fsm_output[0]) | or_tmp_35);
  assign tensor_buf0_val_and_cse = run_wen & (~ (fsm_output[1]));
  assign and_184_cse = run_wen & (~ (fsm_output[0]));
  assign nl_operator_11_false_acc_nl_1 = ({1'b1 , widthIn}) + conv_u2s_11_12(~ Tensor_weight_x_COLUMN_x_lpi_1_dfm_mx0w0);
  assign operator_11_false_acc_nl_1 = nl_operator_11_false_acc_nl_1[11:0];
  assign operator_11_false_acc_itm_11_1 = readslicef_12_1_11(operator_11_false_acc_nl_1);
  assign Tensor_weight_x_COLUMN_equal_tmp = Tensor_weight_x_COLUMN_x_lpi_1_dfm ==
      widthIn;
  assign exitL_exit_Tensor_weight_x_ROW_sva_mx0 = ~((~(exit_Tensor_weight_x_ROW_sva_2_mx0w0
      & Tensor_weight_x_COLUMN_equal_tmp)) & main_stage_0_2);
  assign exit_Tensor_weight_x_ROW_sva_2_mx0w0 = ~((Tensor_weight_x_ROW_y_lpi_1_dfm
      != (operator_9_false_1_acc_tmp[8:0])) | (operator_9_false_1_acc_tmp[9]));
  assign nl_operator_9_false_1_acc_tmp = conv_u2s_9_10(heightIn) + 10'b1111111111;
  assign operator_9_false_1_acc_tmp = nl_operator_9_false_1_acc_tmp[9:0];
  assign nl_Tensor_weight_x_COLUMN_acc_1_nl = Tensor_weight_x_COLUMN_x_lpi_1_dfm
      + 11'b00000000001;
  assign Tensor_weight_x_COLUMN_acc_1_nl = nl_Tensor_weight_x_COLUMN_acc_1_nl[10:0];
  assign Tensor_weight_x_COLUMN_if_2_mux_1_nl = MUX_v_11_2_2(Tensor_weight_x_COLUMN_acc_1_nl,
      ({{10{exit_Tensor_weight_x_ROW_sva_2_mx0w0}}, exit_Tensor_weight_x_ROW_sva_2_mx0w0}),
      Tensor_weight_x_COLUMN_equal_tmp);
  assign Tensor_weight_x_ROW_Tensor_weight_x_ROW_Tensor_weight_x_ROW_Tensor_weight_x_ROW_not_nl
      = ~ exitL_exit_Tensor_weight_x_ROW_sva_mx0;
  assign Tensor_weight_x_COLUMN_x_lpi_1_dfm_mx0w0 = MUX_v_11_2_2(11'b00000000000,
      Tensor_weight_x_COLUMN_if_2_mux_1_nl, Tensor_weight_x_ROW_Tensor_weight_x_ROW_Tensor_weight_x_ROW_Tensor_weight_x_ROW_not_nl);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_34_sva_1 = Tensor_weight_x_COLUMN_if_1_for_61_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[34]);
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1 = ({Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_94_1
      , Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_0}) + conv_s2s_94_95(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg);
  assign Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1 = nl_Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94:0];
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1 = ({Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_94_1
      , Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_0}) + conv_s2s_94_95(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg);
  assign Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1 = nl_Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94:0];
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1 = ({Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_93_0
      , Tensor_weight_x_COLUMN_if_1_acc_16_itm_1_0}) + conv_s2s_94_95(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg);
  assign Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1 = nl_Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94:0];
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1 = conv_s2s_94_95(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg)
      + conv_s2s_94_95({Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg , 1'b0}) + conv_s2s_94_95(Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_93_0);
  assign Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1 = nl_Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94:0];
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1 = conv_s2s_94_95(Tensor_weight_x_COLUMN_if_1_asn_28_itm_1)
      + conv_s2s_94_95({Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg , 1'b0}) +
      conv_s2s_94_95(Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_93_0);
  assign Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1 = nl_Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94:0];
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_68_sva_1 = Tensor_weight_x_COLUMN_if_1_for_27_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[68]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_72_sva_1 = Tensor_weight_x_COLUMN_if_1_for_23_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[72]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_70_sva_1 = Tensor_weight_x_COLUMN_if_1_for_25_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[70]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_51_sva_1 = Tensor_weight_x_COLUMN_if_1_for_44_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[51]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_66_sva_1 = Tensor_weight_x_COLUMN_if_1_for_29_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[66]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_50_sva_1 = Tensor_weight_x_COLUMN_if_1_for_45_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[50]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_67_sva_1 = Tensor_weight_x_COLUMN_if_1_for_28_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[67]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_49_sva_1 = Tensor_weight_x_COLUMN_if_1_for_46_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[49]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_69_sva_1 = Tensor_weight_x_COLUMN_if_1_for_26_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[69]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_48_sva_1 = Tensor_weight_x_COLUMN_if_1_for_47_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[48]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_83_sva_1 = Tensor_weight_x_COLUMN_if_1_for_12_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[83]);
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1 = ({(~ Tensor_weight_x_COLUMN_if_1_for_1_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_2_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_3_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_4_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_5_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_6_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_7_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_8_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_9_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_12_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_13_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_14_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_15_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_16_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_17_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_18_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_19_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_20_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_21_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_22_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_23_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_24_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_25_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_26_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_27_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_28_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_29_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_30_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_31_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_32_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_33_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_34_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_35_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_36_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_37_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_38_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_39_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_40_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_41_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_42_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_43_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_44_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_45_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_46_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_47_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_48_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_49_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_50_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_51_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_52_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_53_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_54_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_55_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_56_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_57_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_58_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_59_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_60_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_61_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_62_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_63_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_64_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_65_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_66_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_67_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_68_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_69_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_70_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_71_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_72_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_73_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_74_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_75_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_76_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_77_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_78_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_79_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_80_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_81_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_82_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_83_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_84_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_85_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_86_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_87_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_88_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_89_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_90_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_91_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_92_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_93_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_94_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)
      , (~ Tensor_weight_x_COLUMN_if_1_for_95_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva)})
      + 95'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
  assign Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1 = nl_Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[94:0];
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_54_sva_1 = Tensor_weight_x_COLUMN_if_1_for_41_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[54]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_82_sva_1 = Tensor_weight_x_COLUMN_if_1_for_13_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[82]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_64_sva_1 = Tensor_weight_x_COLUMN_if_1_for_31_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[64]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_53_sva_1 = Tensor_weight_x_COLUMN_if_1_for_42_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[53]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_65_sva_1 = Tensor_weight_x_COLUMN_if_1_for_30_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[65]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_52_sva_1 = Tensor_weight_x_COLUMN_if_1_for_43_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[52]);
  assign Tensor_weight_x_COLUMN_if_1_and_70_nl = Tensor_weight_x_COLUMN_if_1_for_15_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[80]);
  assign nl_operator_9_false_acc_138_cse_1 = conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_70_nl)
      + conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_84_sva_1);
  assign operator_9_false_acc_138_cse_1 = nl_operator_9_false_acc_138_cse_1[1:0];
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_84_sva_1 = Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[84]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_73_sva_1 = Tensor_weight_x_COLUMN_if_1_for_22_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[73]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_81_sva_1 = Tensor_weight_x_COLUMN_if_1_for_14_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[81]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_32_sva_1 = Tensor_weight_x_COLUMN_if_1_for_63_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[32]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_44_sva_1 = Tensor_weight_x_COLUMN_if_1_for_51_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[44]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_43_sva_1 = Tensor_weight_x_COLUMN_if_1_for_52_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[43]);
  assign Tensor_weight_x_COLUMN_if_1_and_psp_sva_1 = Tensor_weight_x_COLUMN_if_1_for_1_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[94]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_24_sva_1 = Tensor_weight_x_COLUMN_if_1_for_71_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[24]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_45_sva_1 = Tensor_weight_x_COLUMN_if_1_for_50_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[45]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_46_sva_1 = Tensor_weight_x_COLUMN_if_1_for_49_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[46]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_28_sva_1 = Tensor_weight_x_COLUMN_if_1_for_67_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[28]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_41_sva_1 = Tensor_weight_x_COLUMN_if_1_for_54_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[41]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_8_sva_1 = Tensor_weight_x_COLUMN_if_1_for_87_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[8]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_86_sva_1 = Tensor_weight_x_COLUMN_if_1_for_9_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[86]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_76_sva_1 = Tensor_weight_x_COLUMN_if_1_for_19_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[76]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_18_sva_1 = Tensor_weight_x_COLUMN_if_1_for_77_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[18]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_19_sva_1 = Tensor_weight_x_COLUMN_if_1_for_76_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[19]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_35_sva_1 = Tensor_weight_x_COLUMN_if_1_for_60_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[35]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_90_sva_1 = Tensor_weight_x_COLUMN_if_1_for_5_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[90]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_36_sva_1 = Tensor_weight_x_COLUMN_if_1_for_59_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[36]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_22_sva_1 = Tensor_weight_x_COLUMN_if_1_for_73_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[22]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_79_sva_1 = Tensor_weight_x_COLUMN_if_1_for_16_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[79]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_77_sva_1 = Tensor_weight_x_COLUMN_if_1_for_18_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[77]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_85_sva_1 = Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[85]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_75_sva_1 = Tensor_weight_x_COLUMN_if_1_for_20_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[75]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_17_sva_1 = Tensor_weight_x_COLUMN_if_1_for_78_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[17]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_12_sva_1 = Tensor_weight_x_COLUMN_if_1_for_83_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[12]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_21_sva_1 = Tensor_weight_x_COLUMN_if_1_for_74_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[21]);
  assign Tensor_weight_x_COLUMN_if_1_and_65_seb_1 = Tensor_weight_x_COLUMN_if_1_for_81_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[14]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_87_sva_1 = Tensor_weight_x_COLUMN_if_1_for_8_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[87]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_88_sva_1 = Tensor_weight_x_COLUMN_if_1_for_7_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[88]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_42_sva_1 = Tensor_weight_x_COLUMN_if_1_for_53_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[42]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_78_sva_1 = Tensor_weight_x_COLUMN_if_1_for_17_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[78]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_16_sva_1 = Tensor_weight_x_COLUMN_if_1_for_79_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[16]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_10_sva_1 = Tensor_weight_x_COLUMN_if_1_for_85_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[10]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_39_sva_1 = Tensor_weight_x_COLUMN_if_1_for_56_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[39]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_71_sva_1 = Tensor_weight_x_COLUMN_if_1_for_24_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[71]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_74_sva_1 = Tensor_weight_x_COLUMN_if_1_for_21_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[74]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_9_sva_1 = Tensor_weight_x_COLUMN_if_1_for_86_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[9]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_38_sva_1 = Tensor_weight_x_COLUMN_if_1_for_57_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[38]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_20_sva_1 = Tensor_weight_x_COLUMN_if_1_for_75_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[20]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_37_sva_1 = Tensor_weight_x_COLUMN_if_1_for_58_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[37]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_92_sva_1 = Tensor_weight_x_COLUMN_if_1_for_3_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[92]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_33_sva_1 = Tensor_weight_x_COLUMN_if_1_for_62_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[33]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_4_sva_1 = Tensor_weight_x_COLUMN_if_1_for_91_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[4]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_89_sva_1 = Tensor_weight_x_COLUMN_if_1_for_6_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[89]);
  assign Tensor_weight_x_COLUMN_if_1_and_1_psp_sva_1 = Tensor_weight_x_COLUMN_if_1_for_2_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[93]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_26_sva_1 = Tensor_weight_x_COLUMN_if_1_for_69_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[26]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_25_sva_1 = Tensor_weight_x_COLUMN_if_1_for_70_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[25]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_91_sva_1 = Tensor_weight_x_COLUMN_if_1_for_4_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[91]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_57_sva_1 = Tensor_weight_x_COLUMN_if_1_for_38_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[57]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_56_sva_1 = Tensor_weight_x_COLUMN_if_1_for_39_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[56]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_60_sva_1 = Tensor_weight_x_COLUMN_if_1_for_35_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[60]);
  assign Tensor_weight_x_COLUMN_if_1_and_34_seb_1 = Tensor_weight_x_COLUMN_if_1_for_33_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[62]);
  assign Tensor_weight_x_COLUMN_if_1_and_2_psp_58_sva_1 = Tensor_weight_x_COLUMN_if_1_for_37_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[58]);
  assign operator_9_false_asn_221 = Tensor_weight_x_COLUMN_if_1_for_55_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[40]);
  assign or_tmp_3 = main_stage_0_4 & (~ Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_3)
      & (~ operator_11_false_1_slc_operator_11_false_1_acc_11_itm_3) & (fsm_output[1]);
  assign or_tmp_35 = (~ Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_4)
      & (fsm_output[1]);
  assign or_tmp_36 = Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_4
      & (fsm_output[1]);
  assign Tensor_weight_x_COLUMN_if_1_mux_17_cse = MUX_v_9_2_2(Tensor_weight_x_COLUMN_if_1_ac_int_cctor_1_sva_1,
      z_out_2, fsm_output[1]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_shift_rsci_oswt_cse <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_ac_int_cctor_1_sva_1 <= 9'b000000000;
      Tensor_weight_x_COLUMN_if_1_slc_95_64_5_itm_1 <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_slc_95_64_4_itm_1 <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_slc_95_64_3_itm_1 <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_4 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      exitL_exit_Tensor_weight_x_ROW_sva <= 1'b0;
      tensor0_val_2_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_10_itm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor0_val_1_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor0_val_0_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      reg_tensor_y_rsci_oswt_cse <= 1'b0;
      tensor_buf0_val_127_64_lpi_1_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      operator_9_false_acc_97_itm_1 <= 8'b00000000;
      operator_9_false_acc_96_itm_1_7_6 <= 2'b00;
      operator_9_false_acc_108_itm_1 <= 9'b000000000;
      operator_9_false_acc_107_itm_1 <= 9'b000000000;
      operator_9_false_acc_106_itm_1_8_4 <= 5'b00000;
      operator_9_false_acc_106_itm_1_3_0 <= 4'b0000;
      operator_9_false_acc_105_itm_1 <= 9'b000000000;
      operator_9_false_acc_104_itm_1 <= 9'b000000000;
      operator_9_false_acc_103_itm_1 <= 9'b000000000;
      operator_9_false_acc_102_itm_1 <= 9'b000000000;
      operator_9_false_acc_81_itm_1_7_1 <= 7'b0000000;
      operator_9_false_acc_79_itm_1 <= 6'b000000;
      operator_9_false_acc_68_itm_1 <= 6'b000000;
      operator_9_false_acc_71_itm_1 <= 6'b000000;
      operator_9_false_acc_70_itm_1 <= 6'b000000;
      operator_9_false_acc_78_itm_1 <= 7'b0000000;
      operator_9_false_acc_77_itm_1 <= 7'b0000000;
      operator_9_false_acc_76_itm_1_6_1 <= 6'b000000;
      operator_9_false_acc_76_itm_1_0 <= 1'b0;
      operator_9_false_acc_75_itm_1 <= 7'b0000000;
      operator_9_false_acc_74_itm_1_6_5 <= 2'b00;
      operator_9_false_acc_74_itm_1_2_0 <= 3'b000;
      Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm
          <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_for_95_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_psp_sva <= 95'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva <= 95'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_for_93_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_94_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_89_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_90_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_91_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_92_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_81_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_82_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_83_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_84_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_85_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_86_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_87_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_88_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_65_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_66_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_67_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_68_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_69_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_70_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_71_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_72_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_73_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_74_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_75_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_76_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_77_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_78_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_79_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_80_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_1_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_2_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_3_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_4_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_5_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_6_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_7_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_8_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_9_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_12_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_13_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_14_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_15_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_16_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_17_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_18_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_19_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_20_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_21_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_22_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_23_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_24_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_25_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_26_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_27_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_28_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_29_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_30_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_31_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_32_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_33_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_34_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_35_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_36_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_37_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_38_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_39_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_40_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_41_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_42_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_43_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_44_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_45_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_46_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_47_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_48_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_49_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_50_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_51_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_52_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_53_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_54_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_55_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_56_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_57_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_58_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_59_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_60_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_61_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_62_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_63_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_64_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_asn_28_itm_1 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_16_itm_1_0 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_94_1 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_0 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_94_1 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      reg_shift_rsci_oswt_cse <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_ac_int_cctor_1_sva_1 <= 9'b000000000;
      Tensor_weight_x_COLUMN_if_1_slc_95_64_5_itm_1 <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_slc_95_64_4_itm_1 <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_slc_95_64_3_itm_1 <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_4 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      exitL_exit_Tensor_weight_x_ROW_sva <= 1'b0;
      tensor0_val_2_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_10_itm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor0_val_1_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor0_val_0_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      reg_tensor_y_rsci_oswt_cse <= 1'b0;
      tensor_buf0_val_127_64_lpi_1_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      operator_9_false_acc_97_itm_1 <= 8'b00000000;
      operator_9_false_acc_96_itm_1_7_6 <= 2'b00;
      operator_9_false_acc_108_itm_1 <= 9'b000000000;
      operator_9_false_acc_107_itm_1 <= 9'b000000000;
      operator_9_false_acc_106_itm_1_8_4 <= 5'b00000;
      operator_9_false_acc_106_itm_1_3_0 <= 4'b0000;
      operator_9_false_acc_105_itm_1 <= 9'b000000000;
      operator_9_false_acc_104_itm_1 <= 9'b000000000;
      operator_9_false_acc_103_itm_1 <= 9'b000000000;
      operator_9_false_acc_102_itm_1 <= 9'b000000000;
      operator_9_false_acc_81_itm_1_7_1 <= 7'b0000000;
      operator_9_false_acc_79_itm_1 <= 6'b000000;
      operator_9_false_acc_68_itm_1 <= 6'b000000;
      operator_9_false_acc_71_itm_1 <= 6'b000000;
      operator_9_false_acc_70_itm_1 <= 6'b000000;
      operator_9_false_acc_78_itm_1 <= 7'b0000000;
      operator_9_false_acc_77_itm_1 <= 7'b0000000;
      operator_9_false_acc_76_itm_1_6_1 <= 6'b000000;
      operator_9_false_acc_76_itm_1_0 <= 1'b0;
      operator_9_false_acc_75_itm_1 <= 7'b0000000;
      operator_9_false_acc_74_itm_1_6_5 <= 2'b00;
      operator_9_false_acc_74_itm_1_2_0 <= 3'b000;
      Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm
          <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_for_95_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_psp_sva <= 95'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva <= 95'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_for_93_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_94_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_89_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_90_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_91_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_92_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_81_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_82_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_83_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_84_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_85_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_86_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_87_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_88_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_65_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_66_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_67_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_68_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_69_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_70_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_71_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_72_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_73_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_74_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_75_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_76_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_77_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_78_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_79_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_80_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_1_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_2_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_3_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_4_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_5_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_6_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_7_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_8_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_9_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_12_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_13_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_14_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_15_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_16_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_17_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_18_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_19_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_20_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_21_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_22_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_23_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_24_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_25_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_26_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_27_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_28_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_29_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_30_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_31_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_32_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_33_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_34_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_35_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_36_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_37_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_38_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_39_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_40_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_41_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_42_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_43_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_44_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_45_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_46_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_47_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_48_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_49_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_50_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_51_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_52_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_53_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_54_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_55_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_56_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_57_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_58_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_59_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_60_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_61_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_62_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_63_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_for_64_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_asn_28_itm_1 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_16_itm_1_0 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_94_1 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_0 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_94_1 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_shift_rsci_oswt_cse <= ~((((~ main_stage_0_4) | Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_3
          | operator_11_false_1_slc_operator_11_false_1_acc_11_itm_3) & (fsm_output[1]))
          | ((~(Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_4
          & exitL_exit_Tensor_weight_x_ROW_sva)) & (fsm_output[0])));
      Tensor_weight_x_COLUMN_if_1_ac_int_cctor_1_sva_1 <= z_out_2;
      Tensor_weight_x_COLUMN_if_1_slc_95_64_5_itm_1 <= z_out[95:64];
      Tensor_weight_x_COLUMN_if_1_slc_95_64_4_itm_1 <= Tensor_weight_x_COLUMN_if_1_lshift_3_itm[95:64];
      Tensor_weight_x_COLUMN_if_1_slc_95_64_3_itm_1 <= z_out_1[95:64];
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_4 <= MUX_s_1_2_2(operator_11_false_acc_itm_11_1,
          Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_3, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b <= MUX_v_64_2_2(tensor0_val_2_lpi_1_dfm_1,
          Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_9_nl, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b <= MUX_v_64_2_2(Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_10_itm_1,
          Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_11_nl, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b <= MUX_v_64_2_2(tensor_buf0_val_191_128_lpi_1_dfm,
          tensor_buf0_val_127_64_lpi_1_dfm, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b <= MUX_v_64_2_2(tensor_buf0_val_383_320_lpi_1_dfm,
          tensor0_val_3_lpi_1_dfm_1, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b <= MUX_v_64_2_2(tensor0_val_4_lpi_1_dfm_1,
          Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_8_nl, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b <= MUX_v_64_2_2(tensor_buf0_val_127_64_lpi_1_dfm,
          Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_10_itm_1, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b <= MUX_v_64_2_2(tensor0_val_3_lpi_1_dfm_1,
          Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_7_nl, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b <= MUX_v_64_2_2(tensor0_val_1_lpi_1_dfm_1,
          Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_12_nl, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b <= MUX1HOT_v_64_3_2(tensor0_val_0_lpi_1_dfm_1,
          (tensor_y_rsci_idat_mxwt[383:320]), tensor_buf0_val_383_320_lpi_1_dfm,
          {(fsm_output[0]) , or_tmp_35 , or_tmp_36});
      exitL_exit_Tensor_weight_x_ROW_sva <= MUX_s_1_2_2(exitL_exit_Tensor_weight_x_ROW_sva_mx0,
          main_stage_0_4, fsm_output[1]);
      tensor0_val_2_lpi_1_dfm_1 <= MUX1HOT_v_64_3_2(tensor_buf0_val_383_320_lpi_1_dfm,
          (tensor_y_rsci_idat_mxwt[191:128]), tensor_buf0_val_191_128_lpi_1_dfm,
          {(fsm_output[0]) , or_tmp_35 , or_tmp_36});
      Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_10_itm_1 <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          or_nl, nor_nl);
      tensor0_val_1_lpi_1_dfm_1 <= MUX_v_64_2_2(tensor_buf0_val_127_64_lpi_1_dfm,
          (tensor_y_rsci_idat_mxwt[127:64]), or_tmp_35);
      tensor0_val_0_lpi_1_dfm_1 <= MUX1HOT_v_64_3_2(tensor_buf0_val_191_128_lpi_1_dfm,
          (tensor_y_rsci_idat_mxwt[63:0]), Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_10_itm_1,
          {(fsm_output[0]) , or_tmp_35 , or_tmp_36});
      reg_tensor_y_rsci_oswt_cse <= ~((fsm_output[1]) | operator_11_false_acc_itm_11_1);
      tensor_buf0_val_127_64_lpi_1_dfm <= MUX_v_64_2_2(Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_5_nl,
          tensor0_val_4_lpi_1_dfm_1, fsm_output[1]);
      operator_9_false_acc_97_itm_1 <= nl_operator_9_false_acc_97_itm_1[7:0];
      operator_9_false_acc_96_itm_1_7_6 <= nl_operator_9_false_acc_96_itm_1_7_6[1:0];
      operator_9_false_acc_108_itm_1 <= nl_operator_9_false_acc_108_itm_1[8:0];
      operator_9_false_acc_107_itm_1 <= nl_operator_9_false_acc_107_itm_1[8:0];
      operator_9_false_acc_106_itm_1_8_4 <= nl_operator_9_false_acc_106_itm_1_8_4[4:0];
      operator_9_false_acc_106_itm_1_3_0 <= nl_operator_9_false_acc_106_itm_1_3_0[3:0];
      operator_9_false_acc_105_itm_1 <= nl_operator_9_false_acc_105_itm_1[8:0];
      operator_9_false_acc_104_itm_1 <= nl_operator_9_false_acc_104_itm_1[8:0];
      operator_9_false_acc_103_itm_1 <= MUX_v_9_2_2(operator_9_false_acc_nl, operator_9_false_acc_103_nl,
          fsm_output[1]);
      operator_9_false_acc_102_itm_1 <= MUX_v_9_2_2(operator_9_false_acc_118_nl,
          operator_9_false_acc_102_nl, fsm_output[1]);
      operator_9_false_acc_81_itm_1_7_1 <= nl_operator_9_false_acc_81_itm_1_7_1[6:0];
      operator_9_false_acc_79_itm_1 <= nl_operator_9_false_acc_79_itm_1[5:0];
      operator_9_false_acc_68_itm_1 <= nl_operator_9_false_acc_68_itm_1[5:0];
      operator_9_false_acc_71_itm_1 <= nl_operator_9_false_acc_71_itm_1[5:0];
      operator_9_false_acc_70_itm_1 <= nl_operator_9_false_acc_70_itm_1[5:0];
      operator_9_false_acc_78_itm_1 <= nl_operator_9_false_acc_78_itm_1[6:0];
      operator_9_false_acc_77_itm_1 <= nl_operator_9_false_acc_77_itm_1[6:0];
      operator_9_false_acc_76_itm_1_6_1 <= nl_operator_9_false_acc_76_itm_1_6_1[5:0];
      operator_9_false_acc_76_itm_1_0 <= MUX_s_1_2_2((readslicef_11_1_10(operator_11_false_acc_nl)),
          Tensor_weight_x_COLUMN_if_1_and_2_psp_34_sva_1, fsm_output[1]);
      operator_9_false_acc_75_itm_1 <= nl_operator_9_false_acc_75_itm_1[6:0];
      operator_9_false_acc_74_itm_1_6_5 <= nl_operator_9_false_acc_74_itm_1_6_5[1:0];
      operator_9_false_acc_74_itm_1_2_0 <= nl_operator_9_false_acc_74_itm_1_2_0[2:0];
      Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm
          <= MUX_v_32_2_2((readslicef_95_32_63(Tensor_weight_x_COLUMN_if_1_acc_4_nl)),
          Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm_1,
          fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_for_95_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[93]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[93]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[93]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[93]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[93]));
      Tensor_weight_x_COLUMN_if_1_acc_psp_sva <= MUX_v_95_2_2(Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1,
          Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva <= MUX_v_95_2_2(Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1,
          Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_94 <= Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94];
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_93_0 <= MUX_v_94_2_2((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[93:0]),
          Tensor_weight_x_COLUMN_if_1_acc_22_nl, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_94 <= Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94];
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_93_0 <= MUX_v_94_2_2((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[93:0]),
          Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z_oreg, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_94 <= Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94];
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_93_0 <= MUX_v_94_2_2((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[93:0]),
          Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z_oreg, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_for_93_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[91]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[91]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[91]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[91]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[91]));
      Tensor_weight_x_COLUMN_if_1_for_94_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[92]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[92]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[92]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[92]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[92]));
      Tensor_weight_x_COLUMN_if_1_for_89_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[87]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[87]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[87]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[87]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[87]));
      Tensor_weight_x_COLUMN_if_1_for_90_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[88]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[88]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[88]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[88]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[88]));
      Tensor_weight_x_COLUMN_if_1_for_91_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[89]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[89]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[89]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[89]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[89]));
      Tensor_weight_x_COLUMN_if_1_for_92_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[90]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[90]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[90]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[90]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[90]));
      Tensor_weight_x_COLUMN_if_1_for_81_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[79]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[79]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[79]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[79]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[79]));
      Tensor_weight_x_COLUMN_if_1_for_82_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[80]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[80]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[80]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[80]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[80]));
      Tensor_weight_x_COLUMN_if_1_for_83_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[81]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[81]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[81]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[81]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[81]));
      Tensor_weight_x_COLUMN_if_1_for_84_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[82]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[82]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[82]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[82]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[82]));
      Tensor_weight_x_COLUMN_if_1_for_85_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[83]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[83]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[83]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[83]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[83]));
      Tensor_weight_x_COLUMN_if_1_for_86_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[84]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[84]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[84]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[84]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[84]));
      Tensor_weight_x_COLUMN_if_1_for_87_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[85]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[85]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[85]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[85]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[85]));
      Tensor_weight_x_COLUMN_if_1_for_88_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[86]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[86]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[86]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[86]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[86]));
      Tensor_weight_x_COLUMN_if_1_for_65_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[63]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[63]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[63]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[63]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[63]));
      Tensor_weight_x_COLUMN_if_1_for_66_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[64]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[64]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[64]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[64]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[64]));
      Tensor_weight_x_COLUMN_if_1_for_67_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[65]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[65]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[65]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[65]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[65]));
      Tensor_weight_x_COLUMN_if_1_for_68_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[66]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[66]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[66]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[66]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[66]));
      Tensor_weight_x_COLUMN_if_1_for_69_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[67]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[67]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[67]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[67]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[67]));
      Tensor_weight_x_COLUMN_if_1_for_70_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[68]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[68]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[68]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[68]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[68]));
      Tensor_weight_x_COLUMN_if_1_for_71_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[69]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[69]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[69]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[69]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[69]));
      Tensor_weight_x_COLUMN_if_1_for_72_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[70]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[70]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[70]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[70]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[70]));
      Tensor_weight_x_COLUMN_if_1_for_73_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[71]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[71]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[71]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[71]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[71]));
      Tensor_weight_x_COLUMN_if_1_for_74_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[72]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[72]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[72]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[72]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[72]));
      Tensor_weight_x_COLUMN_if_1_for_75_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[73]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[73]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[73]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[73]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[73]));
      Tensor_weight_x_COLUMN_if_1_for_76_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[74]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[74]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[74]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[74]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[74]));
      Tensor_weight_x_COLUMN_if_1_for_77_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[75]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[75]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[75]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[75]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[75]));
      Tensor_weight_x_COLUMN_if_1_for_78_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[76]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[76]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[76]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[76]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[76]));
      Tensor_weight_x_COLUMN_if_1_for_79_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[77]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[77]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[77]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[77]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[77]));
      Tensor_weight_x_COLUMN_if_1_for_80_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[78]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[78]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[78]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[78]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[78]));
      Tensor_weight_x_COLUMN_if_1_for_1_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) | (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94])
          | (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) | (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94])
          | (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]);
      Tensor_weight_x_COLUMN_if_1_for_2_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[0]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[0]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[0]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[0]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[0]));
      Tensor_weight_x_COLUMN_if_1_for_3_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[1]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[1]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[1]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[1]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[1]));
      Tensor_weight_x_COLUMN_if_1_for_4_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[2]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[2]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[2]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[2]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[2]));
      Tensor_weight_x_COLUMN_if_1_for_5_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[3]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[3]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[3]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[3]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[3]));
      Tensor_weight_x_COLUMN_if_1_for_6_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[4]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[4]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[4]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[4]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[4]));
      Tensor_weight_x_COLUMN_if_1_for_7_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[5]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[5]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[5]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[5]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[5]));
      Tensor_weight_x_COLUMN_if_1_for_8_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[6]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[6]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[6]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[6]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[6]));
      Tensor_weight_x_COLUMN_if_1_for_9_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[7]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[7]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[7]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[7]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[7]));
      Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= MUX_s_1_2_2(Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_nl,
          Tensor_weight_x_COLUMN_if_1_and_2_psp_68_sva_1, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= MUX_s_1_2_2(Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_nl,
          Tensor_weight_x_COLUMN_if_1_and_2_psp_72_sva_1, fsm_output[1]);
      Tensor_weight_x_COLUMN_if_1_for_12_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[10]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[10]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[10]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[10]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[10]));
      Tensor_weight_x_COLUMN_if_1_for_13_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[11]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[11]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[11]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[11]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[11]));
      Tensor_weight_x_COLUMN_if_1_for_14_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[12]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[12]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[12]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[12]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[12]));
      Tensor_weight_x_COLUMN_if_1_for_15_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[13]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[13]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[13]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[13]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[13]));
      Tensor_weight_x_COLUMN_if_1_for_16_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[14]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[14]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[14]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[14]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[14]));
      Tensor_weight_x_COLUMN_if_1_for_17_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[15]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[15]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[15]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[15]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[15]));
      Tensor_weight_x_COLUMN_if_1_for_18_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[16]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[16]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[16]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[16]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[16]));
      Tensor_weight_x_COLUMN_if_1_for_19_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[17]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[17]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[17]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[17]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[17]));
      Tensor_weight_x_COLUMN_if_1_for_20_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[18]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[18]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[18]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[18]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[18]));
      Tensor_weight_x_COLUMN_if_1_for_21_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[19]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[19]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[19]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[19]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[19]));
      Tensor_weight_x_COLUMN_if_1_for_22_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[20]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[20]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[20]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[20]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[20]));
      Tensor_weight_x_COLUMN_if_1_for_23_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[21]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[21]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[21]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[21]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[21]));
      Tensor_weight_x_COLUMN_if_1_for_24_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[22]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[22]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[22]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[22]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[22]));
      Tensor_weight_x_COLUMN_if_1_for_25_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[23]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[23]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[23]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[23]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[23]));
      Tensor_weight_x_COLUMN_if_1_for_26_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[24]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[24]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[24]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[24]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[24]));
      Tensor_weight_x_COLUMN_if_1_for_27_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[25]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[25]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[25]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[25]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[25]));
      Tensor_weight_x_COLUMN_if_1_for_28_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[26]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[26]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[26]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[26]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[26]));
      Tensor_weight_x_COLUMN_if_1_for_29_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[27]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[27]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[27]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[27]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[27]));
      Tensor_weight_x_COLUMN_if_1_for_30_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[28]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[28]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[28]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[28]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[28]));
      Tensor_weight_x_COLUMN_if_1_for_31_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[29]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[29]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[29]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[29]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[29]));
      Tensor_weight_x_COLUMN_if_1_for_32_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[30]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[30]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[30]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[30]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[30]));
      Tensor_weight_x_COLUMN_if_1_for_33_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[31]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[31]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[31]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[31]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[31]));
      Tensor_weight_x_COLUMN_if_1_for_34_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[32]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[32]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[32]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[32]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[32]));
      Tensor_weight_x_COLUMN_if_1_for_35_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[33]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[33]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[33]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[33]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[33]));
      Tensor_weight_x_COLUMN_if_1_for_36_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[34]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[34]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[34]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[34]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[34]));
      Tensor_weight_x_COLUMN_if_1_for_37_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[35]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[35]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[35]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[35]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[35]));
      Tensor_weight_x_COLUMN_if_1_for_38_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[36]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[36]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[36]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[36]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[36]));
      Tensor_weight_x_COLUMN_if_1_for_39_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[37]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[37]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[37]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[37]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[37]));
      Tensor_weight_x_COLUMN_if_1_for_40_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[38]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[38]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[38]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[38]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[38]));
      Tensor_weight_x_COLUMN_if_1_for_41_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[39]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[39]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[39]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[39]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[39]));
      Tensor_weight_x_COLUMN_if_1_for_42_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[40]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[40]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[40]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[40]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[40]));
      Tensor_weight_x_COLUMN_if_1_for_43_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[41]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[41]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[41]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[41]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[41]));
      Tensor_weight_x_COLUMN_if_1_for_44_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[42]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[42]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[42]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[42]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[42]));
      Tensor_weight_x_COLUMN_if_1_for_45_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[43]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[43]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[43]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[43]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[43]));
      Tensor_weight_x_COLUMN_if_1_for_46_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[44]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[44]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[44]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[44]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[44]));
      Tensor_weight_x_COLUMN_if_1_for_47_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[45]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[45]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[45]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[45]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[45]));
      Tensor_weight_x_COLUMN_if_1_for_48_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[46]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[46]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[46]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[46]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[46]));
      Tensor_weight_x_COLUMN_if_1_for_49_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[47]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[47]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[47]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[47]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[47]));
      Tensor_weight_x_COLUMN_if_1_for_50_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[48]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[48]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[48]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[48]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[48]));
      Tensor_weight_x_COLUMN_if_1_for_51_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[49]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[49]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[49]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[49]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[49]));
      Tensor_weight_x_COLUMN_if_1_for_52_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[50]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[50]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[50]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[50]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[50]));
      Tensor_weight_x_COLUMN_if_1_for_53_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[51]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[51]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[51]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[51]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[51]));
      Tensor_weight_x_COLUMN_if_1_for_54_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[52]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[52]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[52]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[52]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[52]));
      Tensor_weight_x_COLUMN_if_1_for_55_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[53]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[53]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[53]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[53]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[53]));
      Tensor_weight_x_COLUMN_if_1_for_56_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[54]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[54]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[54]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[54]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[54]));
      Tensor_weight_x_COLUMN_if_1_for_57_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[55]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[55]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[55]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[55]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[55]));
      Tensor_weight_x_COLUMN_if_1_for_58_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[56]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[56]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[56]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[56]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[56]));
      Tensor_weight_x_COLUMN_if_1_for_59_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[57]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[57]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[57]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[57]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[57]));
      Tensor_weight_x_COLUMN_if_1_for_60_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[58]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[58]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[58]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[58]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[58]));
      Tensor_weight_x_COLUMN_if_1_for_61_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[59]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[59]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[59]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[59]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[59]));
      Tensor_weight_x_COLUMN_if_1_for_62_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[60]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[60]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[60]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[60]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[60]));
      Tensor_weight_x_COLUMN_if_1_for_63_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[61]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[61]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[61]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[61]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[61]));
      Tensor_weight_x_COLUMN_if_1_for_64_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
          <= ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[62]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[62]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[62]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[62]))
          | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[62]));
      Tensor_weight_x_COLUMN_if_1_asn_28_itm_1 <= Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z_oreg;
      Tensor_weight_x_COLUMN_if_1_acc_16_itm_1_0 <= Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg[0];
      Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_94_1 <= nl_Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_94_1[93:0];
      Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_0 <= Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg[0];
      Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_94_1 <= nl_Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_94_1[93:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      shift_rsci_idat <= 9'b000000000;
      tensor_shift_rsci_idat_191_160 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_159_128 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_63_32 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_127_96 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_95_64 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      shift_rsci_idat <= 9'b000000000;
      tensor_shift_rsci_idat_191_160 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_159_128 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_63_32 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_127_96 <= 32'b00000000000000000000000000000000;
      tensor_shift_rsci_idat_95_64 <= 32'b00000000000000000000000000000000;
    end
    else if ( Tensor_weight_x_COLUMN_if_1_and_95_cse ) begin
      shift_rsci_idat <= MUX_v_9_2_2(9'b000000000, Tensor_weight_x_COLUMN_if_1_ac_int_cctor_1_sva_1,
          Tensor_weight_x_COLUMN_if_1_not_9_nl);
      tensor_shift_rsci_idat_191_160 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          Tensor_weight_x_COLUMN_if_1_slc_95_64_5_itm_1, Tensor_weight_x_COLUMN_if_1_not_10_nl);
      tensor_shift_rsci_idat_31_0 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (z_out[95:64]), Tensor_weight_x_COLUMN_if_1_not_11_nl);
      tensor_shift_rsci_idat_159_128 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          Tensor_weight_x_COLUMN_if_1_slc_95_64_4_itm_1, Tensor_weight_x_COLUMN_if_1_not_12_nl);
      tensor_shift_rsci_idat_63_32 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (z_out_1[95:64]), Tensor_weight_x_COLUMN_if_1_not_13_nl);
      tensor_shift_rsci_idat_127_96 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          Tensor_weight_x_COLUMN_if_1_slc_95_64_3_itm_1, Tensor_weight_x_COLUMN_if_1_not_14_nl);
      tensor_shift_rsci_idat_95_64 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm,
          Tensor_weight_x_COLUMN_if_1_not_15_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_3 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_2 <= 1'b0;
      tensor_buf1_val_255_192_lpi_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_buf1_val_127_64_lpi_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_buf1_val_63_0_lpi_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_1 <= 1'b0;
      operator_11_false_1_slc_operator_11_false_1_acc_11_itm_3 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm_1
          <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1 <= 95'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1 <= 95'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_0 <= 1'b0;
      operator_11_false_1_slc_operator_11_false_1_acc_11_itm_1 <= 1'b0;
    end
    else if ( rst ) begin
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_3 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_2 <= 1'b0;
      tensor_buf1_val_255_192_lpi_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_buf1_val_127_64_lpi_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_buf1_val_63_0_lpi_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_1 <= 1'b0;
      operator_11_false_1_slc_operator_11_false_1_acc_11_itm_3 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_94 <= 1'b0;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_93_0 <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm_1
          <= 32'b00000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1 <= 95'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1 <= 95'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_0 <= 1'b0;
      operator_11_false_1_slc_operator_11_false_1_acc_11_itm_1 <= 1'b0;
    end
    else if ( Tensor_weight_x_COLUMN_if_1_and_105_cse ) begin
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_3 <= Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_2;
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_2 <= Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_1;
      tensor_buf1_val_255_192_lpi_1 <= tensor0_val_3_lpi_1_dfm_1;
      tensor_buf1_val_127_64_lpi_1 <= tensor_buf0_val_127_64_lpi_1_dfm;
      tensor_buf1_val_63_0_lpi_1 <= Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_10_itm_1;
      Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_1 <= (readslicef_12_1_11(Tensor_weight_x_COLUMN_aelse_acc_nl))
          & (~ operator_9_false_acc_76_itm_1_0);
      operator_11_false_1_slc_operator_11_false_1_acc_11_itm_3 <= Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_0;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_94 <= Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_94;
      Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1_93_0 <= Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_93_0;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_94 <= Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_94;
      Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1_93_0 <= Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_93_0;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_94 <= Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_94;
      Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1_93_0 <= Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_93_0;
      Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm_1
          <= Tensor_weight_x_COLUMN_if_1_slc_Tensor_weight_x_COLUMN_if_1_acc_4_psp_94_63_itm;
      Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1 <= Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva;
      Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1 <= Tensor_weight_x_COLUMN_if_1_acc_psp_sva;
      Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_0 <= MUX_s_1_2_2(operator_11_false_1_slc_operator_11_false_1_acc_11_itm_1,
          (Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg[0]), Tensor_weight_x_COLUMN_if_1_Tensor_weight_x_COLUMN_if_1_and_itm_1);
      operator_11_false_1_slc_operator_11_false_1_acc_11_itm_1 <= readslicef_12_1_11(operator_11_false_1_acc_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      tensor0_val_4_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor0_val_3_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      tensor0_val_4_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor0_val_3_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( tensor0_val_and_cse ) begin
      tensor0_val_4_lpi_1_dfm_1 <= MUX_v_64_2_2(Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_2_nl,
          (tensor_y_rsci_idat_mxwt[319:256]), or_tmp_35);
      tensor0_val_3_lpi_1_dfm_1 <= MUX_v_64_2_2(Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_3_nl,
          (tensor_y_rsci_idat_mxwt[255:192]), or_tmp_35);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      tensor_buf0_val_383_320_lpi_1_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_x_lpi_1_dfm <= 11'b00000000000;
      tensor_buf0_val_191_128_lpi_1_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_ROW_y_lpi_1_dfm <= 9'b000000000;
    end
    else if ( rst ) begin
      tensor_buf0_val_383_320_lpi_1_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_COLUMN_x_lpi_1_dfm <= 11'b00000000000;
      tensor_buf0_val_191_128_lpi_1_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_x_ROW_y_lpi_1_dfm <= 9'b000000000;
    end
    else if ( tensor_buf0_val_and_cse ) begin
      tensor_buf0_val_383_320_lpi_1_dfm <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b, Tensor_weight_x_ROW_not_42_nl);
      Tensor_weight_x_COLUMN_x_lpi_1_dfm <= Tensor_weight_x_COLUMN_x_lpi_1_dfm_mx0w0;
      tensor_buf0_val_191_128_lpi_1_dfm <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          tensor0_val_2_lpi_1_dfm_1, Tensor_weight_x_ROW_not_43_nl);
      Tensor_weight_x_ROW_y_lpi_1_dfm <= MUX_v_9_2_2(9'b000000000, Tensor_weight_x_COLUMN_if_2_mux_nl,
          Tensor_weight_x_ROW_not_34_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
    end
    else if ( rst ) begin
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
    end
    else if ( and_184_cse ) begin
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
    end
  end
  assign Tensor_weight_x_ROW_not_46_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva;
  assign Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_9_nl = MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      tensor_buf1_val_255_192_lpi_1, Tensor_weight_x_ROW_not_46_nl);
  assign Tensor_weight_x_ROW_not_47_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva;
  assign Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_11_nl = MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      tensor_buf1_val_127_64_lpi_1, Tensor_weight_x_ROW_not_47_nl);
  assign Tensor_weight_x_ROW_not_45_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva;
  assign Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_8_nl = MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      tensor0_val_1_lpi_1_dfm_1, Tensor_weight_x_ROW_not_45_nl);
  assign Tensor_weight_x_ROW_not_44_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva;
  assign Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_7_nl = MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      tensor0_val_2_lpi_1_dfm_1, Tensor_weight_x_ROW_not_44_nl);
  assign Tensor_weight_x_ROW_not_48_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva;
  assign Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_12_nl = MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      tensor_buf1_val_63_0_lpi_1, Tensor_weight_x_ROW_not_48_nl);
  assign nor_1_nl = ~(((~ exitL_exit_Tensor_weight_x_ROW_sva) & (fsm_output[1]))
      | ((~ exitL_exit_Tensor_weight_x_ROW_sva_mx0) & (fsm_output[0])));
  assign or_nl = MUX_v_64_2_2(tensor0_val_0_lpi_1_dfm_1, 64'b1111111111111111111111111111111111111111111111111111111111111111,
      nor_1_nl);
  assign nor_nl = ~((exitL_exit_Tensor_weight_x_ROW_sva & (fsm_output[1])) | (exitL_exit_Tensor_weight_x_ROW_sva_mx0
      & (fsm_output[0])));
  assign Tensor_weight_x_ROW_not_40_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva_mx0;
  assign Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_5_nl = MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      tensor0_val_1_lpi_1_dfm_1, Tensor_weight_x_ROW_not_40_nl);
  assign Tensor_weight_x_COLUMN_if_1_and_47_nl = Tensor_weight_x_COLUMN_if_1_for_72_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[23]);
  assign nl_operator_9_false_acc_135_nl = conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_45_sva_1
      , (signext_2_1(Tensor_weight_x_COLUMN_if_1_and_47_nl))}) + conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_46_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_28_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_28_sva_1})});
  assign operator_9_false_acc_135_nl = nl_operator_9_false_acc_135_nl[3:0];
  assign nl_operator_9_false_acc_97_itm_1  = conv_u2u_7_8({operator_9_false_acc_135_nl
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_28_sva_1 , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_28_sva_1})
      + conv_u2u_6_8({Tensor_weight_x_COLUMN_if_1_and_2_psp_43_sva_1 , ({{4{Tensor_weight_x_COLUMN_if_1_and_psp_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_psp_sva_1})}) + conv_u2u_6_8({Tensor_weight_x_COLUMN_if_1_and_2_psp_44_sva_1
      , (signext_5_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_24_sva_1 , 2'b00 , Tensor_weight_x_COLUMN_if_1_and_2_psp_24_sva_1}))});
  assign nl_operator_9_false_acc_96_itm_1_7_6  = conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_68_sva_1)
      + conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_72_sva_1);
  assign nl_operator_9_false_acc_141_nl = conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_73_sva_1)
      + conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_81_sva_1);
  assign operator_9_false_acc_141_nl = nl_operator_9_false_acc_141_nl[1:0];
  assign nl_operator_9_false_acc_142_nl = conv_u2u_2_3({Tensor_weight_x_COLUMN_if_1_and_2_psp_73_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_32_sva_1}) + conv_u2u_2_3({Tensor_weight_x_COLUMN_if_1_and_2_psp_81_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_44_sva_1});
  assign operator_9_false_acc_142_nl = nl_operator_9_false_acc_142_nl[2:0];
  assign nl_operator_9_false_acc_108_itm_1  = conv_u2u_8_9({operator_9_false_acc_138_cse_1
      , operator_9_false_acc_138_cse_1 , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_84_sva_1
      , operator_9_false_acc_138_cse_1}) + conv_u2u_8_9({operator_9_false_acc_141_nl
      , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_81_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_73_sva_1
      , operator_9_false_acc_142_nl});
  assign Tensor_weight_x_COLUMN_if_1_and_36_nl = Tensor_weight_x_COLUMN_if_1_for_32_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[63]);
  assign nl_operator_9_false_acc_143_nl = conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_83_sva_1
      , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_83_sva_1}) + conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_36_nl
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_54_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_54_sva_1})});
  assign operator_9_false_acc_143_nl = nl_operator_9_false_acc_143_nl[3:0];
  assign nl_operator_9_false_acc_144_nl = conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_83_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_82_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_82_sva_1})})
      + conv_u2u_3_4({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_54_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_54_sva_1});
  assign operator_9_false_acc_144_nl = nl_operator_9_false_acc_144_nl[3:0];
  assign nl_operator_9_false_acc_145_nl = conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_64_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_53_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_53_sva_1})})
      + conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_65_sva_1 , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_52_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_52_sva_1})});
  assign operator_9_false_acc_145_nl = nl_operator_9_false_acc_145_nl[3:0];
  assign nl_operator_9_false_acc_146_nl = conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_53_sva_1)
      + conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_52_sva_1);
  assign operator_9_false_acc_146_nl = nl_operator_9_false_acc_146_nl[1:0];
  assign nl_operator_9_false_acc_107_itm_1  = conv_u2u_8_9({operator_9_false_acc_143_nl
      , operator_9_false_acc_144_nl}) + conv_u2u_8_9({operator_9_false_acc_145_nl
      , operator_9_false_acc_146_nl , Tensor_weight_x_COLUMN_if_1_and_2_psp_53_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_52_sva_1});
  assign nl_operator_9_false_acc_106_itm_1_8_4  = conv_u2u_3_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_70_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_51_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_51_sva_1})})
      + conv_u2u_3_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_66_sva_1 , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_50_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_50_sva_1})}) + conv_u2u_3_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_67_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_49_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_49_sva_1})})
      + conv_u2u_3_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_69_sva_1 , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_48_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_48_sva_1})});
  assign nl_operator_9_false_acc_106_itm_1_3_0  = conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_51_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_50_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_50_sva_1})
      + conv_u2u_2_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_49_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_48_sva_1});
  assign Tensor_weight_x_COLUMN_if_1_and_4_nl = Tensor_weight_x_COLUMN_if_1_for_48_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[47]);
  assign nl_operator_9_false_acc_120_nl = conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_71_sva_1
      , (signext_2_1(Tensor_weight_x_COLUMN_if_1_and_4_nl))}) + conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_78_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_34_seb_1}}, Tensor_weight_x_COLUMN_if_1_and_34_seb_1})});
  assign operator_9_false_acc_120_nl = nl_operator_9_false_acc_120_nl[3:0];
  assign Tensor_weight_x_COLUMN_if_1_and_32_nl = Tensor_weight_x_COLUMN_if_1_for_34_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[61]);
  assign nl_operator_9_false_acc_105_itm_1  = conv_u2u_8_9({operator_9_false_acc_120_nl
      , Tensor_weight_x_COLUMN_if_1_and_34_seb_1 , Tensor_weight_x_COLUMN_if_1_and_34_seb_1
      , Tensor_weight_x_COLUMN_if_1_and_34_seb_1 , Tensor_weight_x_COLUMN_if_1_and_34_seb_1})
      + conv_u2u_7_9({Tensor_weight_x_COLUMN_if_1_and_2_psp_74_sva_1 , (signext_6_2({Tensor_weight_x_COLUMN_if_1_and_32_nl
      , 1'b0}))}) + conv_u2u_7_9({Tensor_weight_x_COLUMN_if_1_and_2_psp_77_sva_1
      , (signext_6_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_58_sva_1 , 1'b0 , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_58_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_58_sva_1})}))});
  assign nl_operator_9_false_acc_121_nl = conv_u2u_4_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_75_sva_1
      , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_57_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_57_sva_1})})
      + conv_u2u_4_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_76_sva_1 , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_56_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_56_sva_1})});
  assign operator_9_false_acc_121_nl = nl_operator_9_false_acc_121_nl[4:0];
  assign Tensor_weight_x_COLUMN_if_1_and_20_nl = Tensor_weight_x_COLUMN_if_1_for_40_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[55]);
  assign nl_operator_9_false_acc_122_nl = conv_u2u_4_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_79_sva_1
      , (signext_3_1(Tensor_weight_x_COLUMN_if_1_and_20_nl))}) + conv_u2u_4_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_82_sva_1
      , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_60_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_60_sva_1})});
  assign operator_9_false_acc_122_nl = nl_operator_9_false_acc_122_nl[4:0];
  assign nl_operator_9_false_acc_104_itm_1  = conv_u2u_8_9({operator_9_false_acc_121_nl
      , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_57_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_56_sva_1})
      + conv_u2u_8_9({operator_9_false_acc_122_nl , Tensor_weight_x_COLUMN_if_1_and_2_psp_60_sva_1
      , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_60_sva_1});
  assign nl_operator_9_false_acc_117_nl = z_out_2 + operator_9_false_acc_105_itm_1
      + operator_9_false_acc_104_itm_1;
  assign operator_9_false_acc_117_nl = nl_operator_9_false_acc_117_nl[8:0];
  assign nl_operator_9_false_acc_101_nl = conv_s2s_6_8(operator_9_false_acc_79_itm_1)
      + conv_u2s_6_8(operator_9_false_acc_68_itm_1);
  assign operator_9_false_acc_101_nl = nl_operator_9_false_acc_101_nl[7:0];
  assign nl_operator_9_false_acc_111_nl = conv_u2s_8_9({operator_9_false_acc_81_itm_1_7_1
      , 1'b0}) + conv_s2s_8_9(operator_9_false_acc_101_nl);
  assign operator_9_false_acc_111_nl = nl_operator_9_false_acc_111_nl[8:0];
  assign nl_operator_9_false_acc_100_nl = conv_u2u_7_8(operator_9_false_acc_78_itm_1)
      + conv_u2u_6_8(operator_9_false_acc_71_itm_1) + conv_u2u_6_8(operator_9_false_acc_70_itm_1);
  assign operator_9_false_acc_100_nl = nl_operator_9_false_acc_100_nl[7:0];
  assign nl_operator_9_false_acc_116_nl = operator_9_false_acc_111_nl + conv_u2s_8_9(operator_9_false_acc_100_nl);
  assign operator_9_false_acc_116_nl = nl_operator_9_false_acc_116_nl[8:0];
  assign nl_operator_9_false_acc_110_nl = conv_u2u_7_9(operator_9_false_acc_77_itm_1)
      + conv_u2u_7_9({operator_9_false_acc_76_itm_1_6_1 , operator_9_false_acc_76_itm_1_0})
      + conv_u2u_7_9(operator_9_false_acc_75_itm_1) + conv_u2u_7_9({operator_9_false_acc_74_itm_1_6_5
      , operator_9_false_acc_74_itm_1_6_5 , operator_9_false_acc_74_itm_1_2_0});
  assign operator_9_false_acc_110_nl = nl_operator_9_false_acc_110_nl[8:0];
  assign nl_operator_9_false_acc_119_nl = operator_9_false_acc_116_nl + operator_9_false_acc_110_nl;
  assign operator_9_false_acc_119_nl = nl_operator_9_false_acc_119_nl[8:0];
  assign nl_operator_9_false_acc_nl = operator_9_false_acc_117_nl + operator_9_false_acc_119_nl;
  assign operator_9_false_acc_nl = nl_operator_9_false_acc_nl[8:0];
  assign Tensor_weight_x_COLUMN_if_1_and_28_nl = Tensor_weight_x_COLUMN_if_1_for_36_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[59]);
  assign Tensor_weight_x_COLUMN_if_1_and_31_nl = Tensor_weight_x_COLUMN_if_1_for_64_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[31]);
  assign Tensor_weight_x_COLUMN_if_1_and_39_nl = Tensor_weight_x_COLUMN_if_1_for_68_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[27]);
  assign nl_operator_9_false_acc_123_nl = conv_u2u_5_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_85_sva_1
      , (signext_4_1(Tensor_weight_x_COLUMN_if_1_and_28_nl))}) + conv_u2u_5_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_86_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_31_nl , (signext_3_1(Tensor_weight_x_COLUMN_if_1_and_39_nl))});
  assign operator_9_false_acc_123_nl = nl_operator_9_false_acc_123_nl[5:0];
  assign Tensor_weight_x_COLUMN_if_1_and_33_nl = Tensor_weight_x_COLUMN_if_1_for_65_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[30]);
  assign Tensor_weight_x_COLUMN_if_1_and_35_nl = Tensor_weight_x_COLUMN_if_1_for_66_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[29]);
  assign nl_operator_9_false_acc_103_nl = conv_u2u_8_9({operator_9_false_acc_123_nl
      , 2'b00}) + conv_u2u_7_9({Tensor_weight_x_COLUMN_if_1_and_2_psp_87_sva_1 ,
      Tensor_weight_x_COLUMN_if_1_and_2_psp_32_sva_1 , (signext_5_1(Tensor_weight_x_COLUMN_if_1_and_33_nl))})
      + conv_u2u_7_9({Tensor_weight_x_COLUMN_if_1_and_2_psp_88_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_33_sva_1
      , (signext_5_2({Tensor_weight_x_COLUMN_if_1_and_35_nl , 1'b0}))});
  assign operator_9_false_acc_103_nl = nl_operator_9_false_acc_103_nl[8:0];
  assign nl_operator_9_false_acc_118_nl = operator_9_false_acc_108_itm_1 + operator_9_false_acc_107_itm_1
      + ({operator_9_false_acc_106_itm_1_8_4 , operator_9_false_acc_106_itm_1_3_0})
      + conv_u2u_8_9(operator_9_false_acc_97_itm_1) + conv_u2u_8_9({operator_9_false_acc_96_itm_1_7_6
      , 2'b00 , Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      , Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      , operator_9_false_acc_96_itm_1_7_6});
  assign operator_9_false_acc_118_nl = nl_operator_9_false_acc_118_nl[8:0];
  assign nl_operator_9_false_acc_124_nl = conv_u2u_4_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_89_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_37_sva_1 , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_26_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_26_sva_1})}) + conv_u2u_4_5({Tensor_weight_x_COLUMN_if_1_and_psp_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_34_sva_1 , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_25_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_25_sva_1})});
  assign operator_9_false_acc_124_nl = nl_operator_9_false_acc_124_nl[4:0];
  assign nl_operator_9_false_acc_125_nl = conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_26_sva_1)
      + conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_25_sva_1);
  assign operator_9_false_acc_125_nl = nl_operator_9_false_acc_125_nl[1:0];
  assign Tensor_weight_x_COLUMN_if_1_and_89_nl = Tensor_weight_x_COLUMN_if_1_for_93_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[2]);
  assign nl_operator_9_false_acc_102_nl = conv_u2u_8_9({operator_9_false_acc_124_nl
      , operator_9_false_acc_125_nl , Tensor_weight_x_COLUMN_if_1_and_2_psp_26_sva_1})
      + conv_u2u_7_9({Tensor_weight_x_COLUMN_if_1_and_2_psp_90_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_35_sva_1
      , ({{3{Tensor_weight_x_COLUMN_if_1_and_1_psp_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_1_psp_sva_1})
      , 1'b0}) + conv_u2u_7_9({Tensor_weight_x_COLUMN_if_1_and_2_psp_91_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_38_sva_1
      , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_91_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_91_sva_1})
      , (signext_2_1(Tensor_weight_x_COLUMN_if_1_and_89_nl))});
  assign operator_9_false_acc_102_nl = nl_operator_9_false_acc_102_nl[8:0];
  assign nl_operator_9_false_acc_81_itm_1_7_1  = conv_u2u_6_7({Tensor_weight_x_COLUMN_if_1_and_2_psp_92_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_39_sva_1 , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_92_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_92_sva_1}) , Tensor_weight_x_COLUMN_if_1_and_2_psp_9_sva_1})
      + conv_u2u_6_7({Tensor_weight_x_COLUMN_if_1_and_1_psp_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_42_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_89_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_89_sva_1})
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_4_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_17_sva_1});
  assign nl_operator_9_false_acc_56_nl = conv_u2u_4_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_74_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_69_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_69_sva_1})
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_88_sva_1}) + conv_u2u_2_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_33_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_4_sva_1}) + conv_u2u_2_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_65_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_16_sva_1});
  assign operator_9_false_acc_56_nl = nl_operator_9_false_acc_56_nl[4:0];
  assign nl_operator_9_false_acc_69_nl = conv_u2s_3_5({Tensor_weight_x_COLUMN_if_1_and_2_psp_67_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_66_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_66_sva_1})})
      + conv_s2s_2_5({(~ Tensor_weight_x_COLUMN_if_1_and_2_psp_89_sva_1) , Tensor_weight_x_COLUMN_if_1_and_2_psp_64_sva_1});
  assign operator_9_false_acc_69_nl = nl_operator_9_false_acc_69_nl[4:0];
  assign nl_operator_9_false_acc_79_itm_1  = conv_u2s_5_6(operator_9_false_acc_56_nl)
      + conv_s2s_5_6(operator_9_false_acc_69_nl);
  assign nl_operator_9_false_acc_68_itm_1  = conv_u2u_5_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_20_sva_1
      , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_20_sva_1 , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_20_sva_1})
      + conv_u2u_5_6(signext_5_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_90_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_37_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_37_sva_1})
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_92_sva_1}));
  assign Tensor_weight_x_COLUMN_if_1_and_79_nl = Tensor_weight_x_COLUMN_if_1_for_88_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[7]);
  assign nl_operator_9_false_acc_71_itm_1  = conv_u2u_4_6(signext_4_3({Tensor_weight_x_COLUMN_if_1_and_2_psp_43_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_74_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_74_sva_1})}))
      + conv_u2u_4_6({Tensor_weight_x_COLUMN_if_1_and_79_nl , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_86_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_86_sva_1})}) + conv_u2u_4_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_8_sva_1
      , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_70_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_70_sva_1})})
      + conv_u2u_4_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_9_sva_1 , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_38_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_38_sva_1})});
  assign Tensor_weight_x_COLUMN_if_1_and_83_nl = Tensor_weight_x_COLUMN_if_1_for_90_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[5]);
  assign nl_operator_9_false_acc_127_nl = conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_42_sva_1
      , (signext_2_1(Tensor_weight_x_COLUMN_if_1_and_83_nl))}) + conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_71_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_85_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_85_sva_1})});
  assign operator_9_false_acc_127_nl = nl_operator_9_false_acc_127_nl[3:0];
  assign Tensor_weight_x_COLUMN_if_1_and_81_nl = Tensor_weight_x_COLUMN_if_1_for_89_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[6]);
  assign nl_operator_9_false_acc_70_itm_1  = conv_u2u_5_6({operator_9_false_acc_127_nl
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_76_sva_1}) + conv_u2u_4_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_10_sva_1
      , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_22_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_22_sva_1})})
      + conv_u2u_4_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_39_sva_1 , (signext_3_1(Tensor_weight_x_COLUMN_if_1_and_81_nl))});
  assign Tensor_weight_x_COLUMN_if_1_and_87_nl = Tensor_weight_x_COLUMN_if_1_for_92_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[3]);
  assign Tensor_weight_x_COLUMN_if_1_and_63_nl = Tensor_weight_x_COLUMN_if_1_for_80_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[15]);
  assign nl_operator_9_false_acc_78_itm_1  = conv_u2u_5_7(signext_5_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_87_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_21_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_21_sva_1})
      , 1'b1})) + conv_u2u_5_7(signext_5_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_88_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_87_nl , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_42_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_42_sva_1})})) + conv_u2u_5_7({Tensor_weight_x_COLUMN_if_1_and_63_nl
      , ({{3{Tensor_weight_x_COLUMN_if_1_and_2_psp_78_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_78_sva_1})})
      + conv_u2u_5_7({Tensor_weight_x_COLUMN_if_1_and_2_psp_16_sva_1 , (signext_4_3({Tensor_weight_x_COLUMN_if_1_and_2_psp_44_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_10_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_10_sva_1})}))});
  assign Tensor_weight_x_COLUMN_if_1_and_71_nl = Tensor_weight_x_COLUMN_if_1_for_84_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[11]);
  assign nl_operator_9_false_acc_128_nl = conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_19_sva_1
      , (signext_2_1(Tensor_weight_x_COLUMN_if_1_and_71_nl))}) + conv_u2u_3_4({Tensor_weight_x_COLUMN_if_1_and_2_psp_21_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_65_seb_1}}, Tensor_weight_x_COLUMN_if_1_and_65_seb_1})});
  assign operator_9_false_acc_128_nl = nl_operator_9_false_acc_128_nl[3:0];
  assign nl_operator_9_false_acc_77_itm_1  = conv_u2u_6_7({operator_9_false_acc_128_nl
      , Tensor_weight_x_COLUMN_if_1_and_65_seb_1 , Tensor_weight_x_COLUMN_if_1_and_65_seb_1})
      + conv_u2u_5_7({Tensor_weight_x_COLUMN_if_1_and_2_psp_17_sva_1 , ({{3{Tensor_weight_x_COLUMN_if_1_and_2_psp_46_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_46_sva_1})}) + conv_u2u_5_7({Tensor_weight_x_COLUMN_if_1_and_2_psp_18_sva_1
      , (signext_4_3({Tensor_weight_x_COLUMN_if_1_and_2_psp_12_sva_1 , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_12_sva_1}))});
  assign Tensor_weight_x_COLUMN_if_1_and_67_nl = Tensor_weight_x_COLUMN_if_1_for_82_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[13]);
  assign nl_operator_9_false_acc_76_itm_1_6_1  = conv_u2u_4_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_22_sva_1
      , (signext_3_1(Tensor_weight_x_COLUMN_if_1_and_67_nl))}) + conv_u2u_4_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_79_sva_1
      , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_77_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_77_sva_1})})
      + conv_u2u_4_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_82_sva_1 , ({{2{Tensor_weight_x_COLUMN_if_1_and_2_psp_45_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_45_sva_1})}) + conv_u2u_4_6({Tensor_weight_x_COLUMN_if_1_and_2_psp_85_sva_1
      , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_75_sva_1}}, Tensor_weight_x_COLUMN_if_1_and_2_psp_75_sva_1})
      , Tensor_weight_x_COLUMN_if_1_and_2_psp_34_sva_1});
  assign nl_operator_11_false_acc_nl = conv_u2u_10_11(Tensor_weight_x_COLUMN_x_lpi_1_dfm_mx0w0[10:1])
      + 11'b11111111111;
  assign operator_11_false_acc_nl = nl_operator_11_false_acc_nl[10:0];
  assign Tensor_weight_x_COLUMN_if_1_and_91_nl = Tensor_weight_x_COLUMN_if_1_for_94_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[1]);
  assign Tensor_weight_x_COLUMN_if_1_and_93_nl = Tensor_weight_x_COLUMN_if_1_for_95_Tensor_weight_x_COLUMN_if_1_for_or_1_psp_sva
      & (Tensor_weight_x_COLUMN_if_1_acc_13_sdt_sva_1[0]);
  assign nl_operator_9_false_acc_75_itm_1  = conv_u2u_6_7({Tensor_weight_x_COLUMN_if_1_and_2_psp_36_sva_1
      , 2'b00 , Tensor_weight_x_COLUMN_if_1_and_2_psp_36_sva_1 , 1'b0 , Tensor_weight_x_COLUMN_if_1_and_2_psp_36_sva_1})
      + conv_u2u_5_7({Tensor_weight_x_COLUMN_if_1_and_2_psp_86_sva_1 , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_76_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_76_sva_1}) , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_18_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_18_sva_1})}) + conv_u2u_3_7({Tensor_weight_x_COLUMN_if_1_and_2_psp_19_sva_1
      , Tensor_weight_x_COLUMN_if_1_and_91_nl , Tensor_weight_x_COLUMN_if_1_and_93_nl})
      + conv_u2u_3_7({Tensor_weight_x_COLUMN_if_1_and_2_psp_35_sva_1 , ({{1{Tensor_weight_x_COLUMN_if_1_and_2_psp_90_sva_1}},
      Tensor_weight_x_COLUMN_if_1_and_2_psp_90_sva_1})});
  assign nl_operator_9_false_acc_74_itm_1_6_5  = conv_u2u_1_2(operator_9_false_asn_221)
      + conv_u2u_1_2(Tensor_weight_x_COLUMN_if_1_and_2_psp_41_sva_1);
  assign nl_operator_9_false_acc_74_itm_1_2_0  = conv_u2u_1_3(operator_9_false_asn_221)
      + conv_u2u_2_3({Tensor_weight_x_COLUMN_if_1_and_2_psp_41_sva_1 , Tensor_weight_x_COLUMN_if_1_and_2_psp_8_sva_1});
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_4_nl = conv_s2s_94_95(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg)
      + conv_s2s_94_95({Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg , 1'b0}) +
      conv_s2s_94_95(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg);
  assign Tensor_weight_x_COLUMN_if_1_acc_4_nl = nl_Tensor_weight_x_COLUMN_if_1_acc_4_nl[94:0];
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_22_nl = conv_s2u_93_94(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z_oreg)
      + conv_s2u_93_94(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z_oreg[93:1]);
  assign Tensor_weight_x_COLUMN_if_1_acc_22_nl = nl_Tensor_weight_x_COLUMN_if_1_acc_22_nl[93:0];
  assign Tensor_weight_x_COLUMN_if_1_for_10_Tensor_weight_x_COLUMN_if_1_for_or_1_nl
      = ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[8]))
      | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[8]))
      | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[8]))
      | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[8]))
      | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[8]));
  assign Tensor_weight_x_COLUMN_if_1_for_11_Tensor_weight_x_COLUMN_if_1_for_or_1_nl
      = ((Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_psp_sva_1_1[9]))
      | ((Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_2_psp_sva_1_1[9]))
      | ((Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_6_psp_sva_1[9]))
      | ((Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_8_psp_sva_1[9]))
      | ((Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[94]) ^ (Tensor_weight_x_COLUMN_if_1_acc_10_psp_sva_1[9]));
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_15_itm_1_94_1  = conv_s2u_93_94(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z_oreg)
      + conv_s2u_93_94(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z_oreg[93:1]);
  assign nl_Tensor_weight_x_COLUMN_if_1_acc_14_itm_1_94_1  = conv_s2u_93_94(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z_oreg)
      + conv_s2u_93_94(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z_oreg[93:1]);
  assign Tensor_weight_x_COLUMN_if_1_not_9_nl = ~ or_tmp_3;
  assign Tensor_weight_x_COLUMN_if_1_not_10_nl = ~ or_tmp_3;
  assign Tensor_weight_x_COLUMN_if_1_not_11_nl = ~ or_tmp_3;
  assign Tensor_weight_x_COLUMN_if_1_not_12_nl = ~ or_tmp_3;
  assign Tensor_weight_x_COLUMN_if_1_not_13_nl = ~ or_tmp_3;
  assign Tensor_weight_x_COLUMN_if_1_not_14_nl = ~ or_tmp_3;
  assign Tensor_weight_x_COLUMN_if_1_not_15_nl = ~ or_tmp_3;
  assign nl_Tensor_weight_x_COLUMN_aelse_acc_nl = ({1'b1 , Tensor_weight_x_COLUMN_x_lpi_1_dfm})
      + conv_u2u_11_12(~ widthIn) + 12'b000000000001;
  assign Tensor_weight_x_COLUMN_aelse_acc_nl = nl_Tensor_weight_x_COLUMN_aelse_acc_nl[11:0];
  assign nl_operator_11_false_1_acc_nl = conv_u2s_11_12(Tensor_weight_x_COLUMN_x_lpi_1_dfm)
      + 12'b111111111111;
  assign operator_11_false_1_acc_nl = nl_operator_11_false_1_acc_nl[11:0];
  assign Tensor_weight_x_ROW_not_38_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva_mx0;
  assign Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_2_nl = MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      tensor0_val_4_lpi_1_dfm_1, Tensor_weight_x_ROW_not_38_nl);
  assign Tensor_weight_x_ROW_not_41_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva_mx0;
  assign Tensor_weight_x_ROW_Tensor_weight_x_ROW_and_3_nl = MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      tensor0_val_3_lpi_1_dfm_1, Tensor_weight_x_ROW_not_41_nl);
  assign Tensor_weight_x_ROW_not_42_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva_mx0;
  assign Tensor_weight_x_ROW_not_43_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva_mx0;
  assign nl_Tensor_weight_x_ROW_acc_nl = Tensor_weight_x_ROW_y_lpi_1_dfm + 9'b000000001;
  assign Tensor_weight_x_ROW_acc_nl = nl_Tensor_weight_x_ROW_acc_nl[8:0];
  assign Tensor_weight_x_COLUMN_if_2_mux_nl = MUX_v_9_2_2(Tensor_weight_x_ROW_y_lpi_1_dfm,
      Tensor_weight_x_ROW_acc_nl, Tensor_weight_x_COLUMN_equal_tmp);
  assign Tensor_weight_x_ROW_not_34_nl = ~ exitL_exit_Tensor_weight_x_ROW_sva_mx0;
  assign nl_z_out_2 = operator_9_false_acc_103_itm_1 + operator_9_false_acc_102_itm_1;
  assign z_out_2 = nl_z_out_2[8:0];

  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | (input_1 & {64{sel[1]}});
    result = result | (input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [93:0] MUX_v_94_2_2;
    input [93:0] input_0;
    input [93:0] input_1;
    input  sel;
    reg [93:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_94_2_2 = result;
  end
  endfunction


  function automatic [94:0] MUX_v_95_2_2;
    input [94:0] input_0;
    input [94:0] input_1;
    input  sel;
    reg [94:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_95_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction


  function automatic [31:0] readslicef_95_32_63;
    input [94:0] vector;
    reg [94:0] tmp;
  begin
    tmp = vector >> 63;
    readslicef_95_32_63 = tmp[31:0];
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input  vector;
  begin
    signext_3_1= {{2{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input  vector;
  begin
    signext_4_1= {{3{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_3;
    input [2:0] vector;
  begin
    signext_4_3= {{1{vector[2]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input  vector;
  begin
    signext_5_1= {{4{vector}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_2;
    input [1:0] vector;
  begin
    signext_5_2= {{3{vector[1]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_4;
    input [3:0] vector;
  begin
    signext_5_4= {{1{vector[3]}}, vector};
  end
  endfunction


  function automatic [5:0] signext_6_2;
    input [1:0] vector;
  begin
    signext_6_2= {{4{vector[1]}}, vector};
  end
  endfunction


  function automatic [5:0] signext_6_4;
    input [3:0] vector;
  begin
    signext_6_4= {{2{vector[3]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2s_2_5 ;
    input [1:0]  vector ;
  begin
    conv_s2s_2_5 = {{3{vector[1]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [7:0] conv_s2s_6_8 ;
    input [5:0]  vector ;
  begin
    conv_s2s_6_8 = {{2{vector[5]}}, vector};
  end
  endfunction


  function automatic [8:0] conv_s2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_9 = {vector[7], vector};
  end
  endfunction


  function automatic [94:0] conv_s2s_94_95 ;
    input [93:0]  vector ;
  begin
    conv_s2s_94_95 = {vector[93], vector};
  end
  endfunction


  function automatic [93:0] conv_s2u_93_94 ;
    input [92:0]  vector ;
  begin
    conv_s2u_93_94 = {vector[92], vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_3_5 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_5 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [5:0] conv_u2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_6 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_6_8 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_8 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_2_5 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_5 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_3_5 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_5 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_3_7 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_7 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_4_6 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_6 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_7 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_6_8 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_8 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_7_9 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_9 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x_struct
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x_struct (
  clk, rst, arst_n, tensor_y_rsc_dat_val, tensor_y_rsc_vld, tensor_y_rsc_rdy, tensor_shift_rsc_dat_val,
      tensor_shift_rsc_vld, tensor_shift_rsc_rdy, shift_rsc_dat, shift_rsc_vld, shift_rsc_rdy,
      widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [383:0] tensor_y_rsc_dat_val;
  input tensor_y_rsc_vld;
  output tensor_y_rsc_rdy;
  output [191:0] tensor_shift_rsc_dat_val;
  output tensor_shift_rsc_vld;
  input tensor_shift_rsc_rdy;
  output [8:0] shift_rsc_dat;
  output shift_rsc_vld;
  input shift_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;


  // Interconnect Declarations
  wire [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b;
  wire [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b;
  wire [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b;
  wire [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b;
  wire [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b;
  wire [63:0] Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b;
  wire [63:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b;
  wire [63:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b;
  wire [63:0] Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b;
  wire [191:0] tensor_shift_rsc_dat;


  // Interconnect Declarations for Component Instantiations 
  wire [94:0] nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z;
  assign nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b);
  wire [94:0] nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z;
  assign nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b);
  wire [94:0] nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z;
  assign nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b);
  wire [94:0] nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z;
  assign nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b);
  wire [94:0] nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z;
  assign nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b);
  wire [94:0] nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z;
  assign nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b);
  wire [93:0] nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z;
  assign nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z
      = $signed(30'b010110011110111011001011111111) * $signed(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b);
  wire [93:0] nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z;
  assign nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z
      = $signed(30'b010110011110111011001011111111) * $signed(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b);
  wire [93:0] nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z;
  assign nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z
      = $signed(30'b010110011110111011001011111111) * $signed(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b);
  OpticalFlow_tensor_weight_x_run OpticalFlow_tensor_weight_x_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_y_rsc_dat(tensor_y_rsc_dat_val),
      .tensor_y_rsc_vld(tensor_y_rsc_vld),
      .tensor_y_rsc_rdy(tensor_y_rsc_rdy),
      .tensor_shift_rsc_dat(tensor_shift_rsc_dat),
      .tensor_shift_rsc_vld(tensor_shift_rsc_vld),
      .tensor_shift_rsc_rdy(tensor_shift_rsc_rdy),
      .shift_rsc_dat(shift_rsc_dat),
      .shift_rsc_vld(shift_rsc_vld),
      .shift_rsc_rdy(shift_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_b),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z(nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_z[93:0]),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_b),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z(nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_1_z[93:0]),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_b),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z(nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_2_z[93:0]),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_b),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z(nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_3_z[93:0]),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_b),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z(nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_4_z[93:0]),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b(Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_b),
      .Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z(nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_2_cmp_5_z[93:0]),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_b),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z(nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_1_cmp_z[92:0]),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_b),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z(nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_1_cmp_1_z[92:0]),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b(Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_b),
      .Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z(nl_OpticalFlow_tensor_weight_x_run_inst_Tensor_weight_x_COLUMN_if_1_mul_1_cmp_2_z[92:0])
    );
  assign tensor_shift_rsc_dat_val = tensor_shift_rsc_dat;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_x
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_x (
  clk, rst, arst_n, tensor_y_rsc_dat, tensor_y_rsc_vld, tensor_y_rsc_rdy, tensor_shift_rsc_dat,
      tensor_shift_rsc_vld, tensor_shift_rsc_rdy, shift_rsc_dat, shift_rsc_vld, shift_rsc_rdy,
      widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [383:0] tensor_y_rsc_dat;
  input tensor_y_rsc_vld;
  output tensor_y_rsc_rdy;
  output [191:0] tensor_shift_rsc_dat;
  output tensor_shift_rsc_vld;
  input tensor_shift_rsc_rdy;
  output [8:0] shift_rsc_dat;
  output shift_rsc_vld;
  input shift_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;


  // Interconnect Declarations
  wire [191:0] tensor_shift_rsc_dat_val;


  // Interconnect Declarations for Component Instantiations 
  OpticalFlow_tensor_weight_x_struct OpticalFlow_tensor_weight_x_struct_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_y_rsc_dat_val(tensor_y_rsc_dat),
      .tensor_y_rsc_vld(tensor_y_rsc_vld),
      .tensor_y_rsc_rdy(tensor_y_rsc_rdy),
      .tensor_shift_rsc_dat_val(tensor_shift_rsc_dat_val),
      .tensor_shift_rsc_vld(tensor_shift_rsc_vld),
      .tensor_shift_rsc_rdy(tensor_shift_rsc_rdy),
      .shift_rsc_dat(shift_rsc_dat),
      .shift_rsc_vld(shift_rsc_vld),
      .shift_rsc_rdy(shift_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn)
    );
  assign tensor_shift_rsc_dat = tensor_shift_rsc_dat_val;
endmodule




//------> ../OpticalFlow_tensor_weight_y.v3/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Mon Jun 17 23:38:03 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_6_9_768_512_1_512_768_1_gen
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_6_9_768_512_1_512_768_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [767:0] q;
  output we;
  output [767:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [767:0] d_d;
  output [767:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_5_9_768_512_1_512_768_1_gen
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_5_9_768_512_1_512_768_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [767:0] q;
  output we;
  output [767:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [767:0] d_d;
  output [767:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for OpticalFlow_tensor_weight_y_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : OpticalFlow_tensor_weight_y_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_run_staller
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_run_staller (
  run_wen, out_product_rsci_wen_comp, tensor_y_rsci_wen_comp
);
  output run_wen;
  input out_product_rsci_wen_comp;
  input tensor_y_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = out_product_rsci_wen_comp & tensor_y_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_run_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_run_wait_dp (
  clk, rst, arst_n, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z, run_wen, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg
);
  input clk;
  input rst;
  input arst_n;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z;
  input run_wen;
  output [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg;
  reg [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg;
  output [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg;
  reg [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg;
  output [92:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg;
  output [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg;
  reg [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg;
  output [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg;
  reg [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg;
  output [92:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg;
  output [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg;
  reg [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg;
  output [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg;
  reg [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg;
  output [92:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg;


  // Interconnect Declarations
  reg [92:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg_pconst_92_0;
  reg [92:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg_pconst_92_0;
  reg [92:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg_pconst_92_0;


  // Interconnect Declarations for Component Instantiations 
  assign Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg = Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg_pconst_92_0;
  assign Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg = Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg_pconst_92_0;
  assign Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg = Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg_pconst_92_0;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg_pconst_92_0 <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg_pconst_92_0 <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg_pconst_92_0 <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg_pconst_92_0 <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg_pconst_92_0 <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg <= 94'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg_pconst_92_0 <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg <= Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg <= Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg_pconst_92_0 <= Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z[92:0];
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg <= Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg <= Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg_pconst_92_0 <= Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z[92:0];
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg <= Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg <= Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg_pconst_92_0 <= Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z[92:0];
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_run_tensor_y_rsci_tensor_y_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_run_tensor_y_rsci_tensor_y_wait_dp (
  clk, rst, arst_n, tensor_y_rsci_oswt, tensor_y_rsci_wen_comp, tensor_y_rsci_biwt,
      tensor_y_rsci_bdwt, tensor_y_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input tensor_y_rsci_oswt;
  output tensor_y_rsci_wen_comp;
  input tensor_y_rsci_biwt;
  input tensor_y_rsci_bdwt;
  output tensor_y_rsci_bcwt;
  reg tensor_y_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign tensor_y_rsci_wen_comp = (~ tensor_y_rsci_oswt) | tensor_y_rsci_biwt | tensor_y_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      tensor_y_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      tensor_y_rsci_bcwt <= 1'b0;
    end
    else begin
      tensor_y_rsci_bcwt <= ~((~(tensor_y_rsci_bcwt | tensor_y_rsci_biwt)) | tensor_y_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_run_tensor_y_rsci_tensor_y_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_run_tensor_y_rsci_tensor_y_wait_ctrl (
  run_wen, tensor_y_rsci_oswt, tensor_y_rsci_biwt, tensor_y_rsci_bdwt, tensor_y_rsci_bcwt,
      tensor_y_rsci_irdy, tensor_y_rsci_ivld_run_sct
);
  input run_wen;
  input tensor_y_rsci_oswt;
  output tensor_y_rsci_biwt;
  output tensor_y_rsci_bdwt;
  input tensor_y_rsci_bcwt;
  input tensor_y_rsci_irdy;
  output tensor_y_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire tensor_y_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign tensor_y_rsci_bdwt = tensor_y_rsci_oswt & run_wen;
  assign tensor_y_rsci_biwt = tensor_y_rsci_ogwt & tensor_y_rsci_irdy;
  assign tensor_y_rsci_ogwt = tensor_y_rsci_oswt & (~ tensor_y_rsci_bcwt);
  assign tensor_y_rsci_ivld_run_sct = tensor_y_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_run_out_product_rsci_out_product_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_run_out_product_rsci_out_product_wait_ctrl (
  run_wen, out_product_rsci_iswt0, out_product_rsci_irdy_run_sct
);
  input run_wen;
  input out_product_rsci_iswt0;
  output out_product_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign out_product_rsci_irdy_run_sct = out_product_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_run_tensor_y_rsci
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_run_tensor_y_rsci (
  clk, rst, arst_n, tensor_y_rsc_dat, tensor_y_rsc_vld, tensor_y_rsc_rdy, run_wen,
      tensor_y_rsci_oswt, tensor_y_rsci_wen_comp, tensor_y_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [383:0] tensor_y_rsc_dat;
  output tensor_y_rsc_vld;
  input tensor_y_rsc_rdy;
  input run_wen;
  input tensor_y_rsci_oswt;
  output tensor_y_rsci_wen_comp;
  input [383:0] tensor_y_rsci_idat;


  // Interconnect Declarations
  wire tensor_y_rsci_biwt;
  wire tensor_y_rsci_bdwt;
  wire tensor_y_rsci_bcwt;
  wire tensor_y_rsci_irdy;
  wire tensor_y_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd384)) tensor_y_rsci (
      .irdy(tensor_y_rsci_irdy),
      .ivld(tensor_y_rsci_ivld_run_sct),
      .idat(tensor_y_rsci_idat),
      .rdy(tensor_y_rsc_rdy),
      .vld(tensor_y_rsc_vld),
      .dat(tensor_y_rsc_dat)
    );
  OpticalFlow_tensor_weight_y_run_tensor_y_rsci_tensor_y_wait_ctrl OpticalFlow_tensor_weight_y_run_tensor_y_rsci_tensor_y_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .tensor_y_rsci_oswt(tensor_y_rsci_oswt),
      .tensor_y_rsci_biwt(tensor_y_rsci_biwt),
      .tensor_y_rsci_bdwt(tensor_y_rsci_bdwt),
      .tensor_y_rsci_bcwt(tensor_y_rsci_bcwt),
      .tensor_y_rsci_irdy(tensor_y_rsci_irdy),
      .tensor_y_rsci_ivld_run_sct(tensor_y_rsci_ivld_run_sct)
    );
  OpticalFlow_tensor_weight_y_run_tensor_y_rsci_tensor_y_wait_dp OpticalFlow_tensor_weight_y_run_tensor_y_rsci_tensor_y_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_y_rsci_oswt(tensor_y_rsci_oswt),
      .tensor_y_rsci_wen_comp(tensor_y_rsci_wen_comp),
      .tensor_y_rsci_biwt(tensor_y_rsci_biwt),
      .tensor_y_rsci_bdwt(tensor_y_rsci_bdwt),
      .tensor_y_rsci_bcwt(tensor_y_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_run_out_product_rsci
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_run_out_product_rsci (
  out_product_rsc_dat, out_product_rsc_vld, out_product_rsc_rdy, run_wen, out_product_rsci_oswt,
      out_product_rsci_wen_comp, out_product_rsci_idat_mxwt
);
  input [383:0] out_product_rsc_dat;
  input out_product_rsc_vld;
  output out_product_rsc_rdy;
  input run_wen;
  input out_product_rsci_oswt;
  output out_product_rsci_wen_comp;
  output [383:0] out_product_rsci_idat_mxwt;


  // Interconnect Declarations
  wire out_product_rsci_irdy_run_sct;
  wire out_product_rsci_ivld;
  wire [383:0] out_product_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd1),
  .width(32'sd384)) out_product_rsci (
      .rdy(out_product_rsc_rdy),
      .vld(out_product_rsc_vld),
      .dat(out_product_rsc_dat),
      .irdy(out_product_rsci_irdy_run_sct),
      .ivld(out_product_rsci_ivld),
      .idat(out_product_rsci_idat)
    );
  OpticalFlow_tensor_weight_y_run_out_product_rsci_out_product_wait_ctrl OpticalFlow_tensor_weight_y_run_out_product_rsci_out_product_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .out_product_rsci_iswt0(out_product_rsci_oswt),
      .out_product_rsci_irdy_run_sct(out_product_rsci_irdy_run_sct)
    );
  assign out_product_rsci_idat_mxwt = out_product_rsci_idat;
  assign out_product_rsci_wen_comp = (~ out_product_rsci_oswt) | out_product_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_run
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_run (
  clk, rst, arst_n, out_product_rsc_dat, out_product_rsc_vld, out_product_rsc_rdy,
      tensor_y_rsc_dat, tensor_y_rsc_vld, tensor_y_rsc_rdy, widthIn, heightIn, line_buf1_rsci_adr_d,
      line_buf1_rsci_clken_d, line_buf1_rsci_d_d, line_buf1_rsci_q_d, line_buf0_rsci_adr_d,
      line_buf0_rsci_d_d, line_buf0_rsci_q_d, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z, Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b,
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z, line_buf1_rsci_we_d_pff, line_buf1_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff,
      line_buf0_rsci_we_d_pff
);
  input clk;
  input rst;
  input arst_n;
  input [383:0] out_product_rsc_dat;
  input out_product_rsc_vld;
  output out_product_rsc_rdy;
  output [383:0] tensor_y_rsc_dat;
  output tensor_y_rsc_vld;
  input tensor_y_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  output [8:0] line_buf1_rsci_adr_d;
  output line_buf1_rsci_clken_d;
  output [767:0] line_buf1_rsci_d_d;
  input [767:0] line_buf1_rsci_q_d;
  output [8:0] line_buf0_rsci_adr_d;
  output [767:0] line_buf0_rsci_d_d;
  input [767:0] line_buf0_rsci_q_d;
  output [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z;
  output [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z;
  output [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z;
  output [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z;
  output [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z;
  output [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z;
  output [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z;
  output [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z;
  output [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b;
  input [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z;
  output line_buf1_rsci_we_d_pff;
  output line_buf1_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff;
  output line_buf0_rsci_we_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire out_product_rsci_wen_comp;
  wire [383:0] out_product_rsci_idat_mxwt;
  wire tensor_y_rsci_wen_comp;
  wire [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg;
  wire [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg;
  wire [92:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg;
  wire [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg;
  wire [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg;
  wire [92:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg;
  wire [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg;
  wire [93:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg;
  wire [92:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg;
  reg [63:0] tensor_y_rsci_idat_383_320;
  reg [63:0] tensor_y_rsci_idat_319_256;
  reg [63:0] tensor_y_rsci_idat_255_192;
  reg [63:0] tensor_y_rsci_idat_191_128;
  reg [63:0] tensor_y_rsci_idat_127_64;
  reg [63:0] tensor_y_rsci_idat_63_0;
  wire [2:0] fsm_output;
  wire Tensor_weight_y_ROW_equal_1_tmp;
  wire Tensor_weight_y_COLUMN_if_4_mux_1_tmp_0;
  wire and_40_cse;
  reg [10:0] Tensor_weight_y_COLUMN_x_lpi_1_dfm;
  wire [11:0] operator_11_false_acc_psp_sva_1;
  wire [12:0] nl_operator_11_false_acc_psp_sva_1;
  wire exitL_exit_Tensor_weight_y_ROW_sva_mx0;
  reg Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1;
  reg operator_9_false_slc_operator_9_false_acc_8_svs_1;
  reg main_stage_0_2;
  reg operator_9_false_slc_operator_9_false_acc_8_svs;
  reg operator_9_false_1_slc_operator_9_false_1_acc_9_itm;
  reg Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_and_itm_1;
  reg main_stage_0_3;
  reg Tensor_weight_y_COLUMN_if_slc_Tensor_weight_y_COLUMN_acc_9_svs;
  reg Tensor_weight_y_COLUMN_x_lpi_1_dfm_1_0;
  wire [8:0] Tensor_weight_y_ROW_y_lpi_1_dfm_mx0w0;
  reg [8:0] Tensor_weight_y_ROW_y_lpi_1_dfm;
  reg [10:0] Tensor_weight_y_COLUMN_x_sva_2_1;
  wire [11:0] nl_Tensor_weight_y_COLUMN_x_sva_2_1;
  wire Tensor_weight_y_COLUMN_if_3_and_cse;
  reg reg_tensor_y_rsci_iswt0_cse;
  reg reg_out_product_rsci_iswt0_cse;
  wire rdbuf0_and_cse;
  wire and_37_cse;
  wire Tensor_weight_y_COLUMN_if_3_and_6_cse;
  wire Tensor_weight_y_COLUMN_qelse_1_and_cse;
  reg [383:0] out_product0_val_lpi_1;
  wire [383:0] out_product0_val_lpi_1_dfm_mx1;
  reg [63:0] wrbuf0_383_320_lpi_1_dfm_2;
  reg [63:0] wrbuf0_319_256_lpi_1_dfm_2;
  reg [63:0] wrbuf0_255_192_lpi_1_dfm_2;
  reg [63:0] wrbuf0_191_128_lpi_1_dfm_2;
  reg [63:0] wrbuf0_127_64_lpi_1_dfm_2;
  reg [63:0] wrbuf0_63_0_lpi_1_dfm_2;
  wire [10:0] Tensor_weight_y_COLUMN_x_lpi_1_dfm_2;
  reg [767:0] rdbuf0_lpi_1;
  wire Tensor_weight_y_COLUMN_if_3_or_itm;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_slc_94_31_5_itm;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_slc_94_31_4_itm;
  reg [63:0] Tensor_weight_y_COLUMN_if_3_slc_94_31_3_itm;
  reg [383:0] out_product0_val_lpi_1_dfm_1;
  reg [383:0] rdbuf1_lpi_1_767_384;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_9_93_30;
  wire [64:0] nl_Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_9_93_30;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_11_93_30;
  wire [64:0] nl_Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_11_93_30;
  reg [191:0] Tensor_weight_y_COLUMN_qr_lpi_1_dfm_383_192;
  reg [191:0] Tensor_weight_y_COLUMN_qr_lpi_1_dfm_191_0;
  reg [191:0] Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_383_192;
  reg [191:0] Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_191_0;
  wire [191:0] Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_mx1_383_192;
  wire [191:0] Tensor_weight_y_COLUMN_qr_lpi_1_dfm_mx1_383_192;
  wire operator_9_false_acc_itm_9_1;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_acc_39_itm_94_31_1;
  wire [63:0] z_out_94_31;
  wire [63:0] z_out_1_94_31;

  wire Tensor_weight_y_COLUMN_if_3_not_6_nl;
  wire Tensor_weight_y_COLUMN_if_3_not_7_nl;
  wire Tensor_weight_y_COLUMN_if_3_not_8_nl;
  wire Tensor_weight_y_COLUMN_if_3_not_9_nl;
  wire Tensor_weight_y_COLUMN_if_3_not_10_nl;
  wire Tensor_weight_y_COLUMN_if_3_not_11_nl;
  wire and_122_nl;
  wire Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_and_nl;
  wire[9:0] Tensor_weight_y_COLUMN_aelse_acc_nl;
  wire[10:0] nl_Tensor_weight_y_COLUMN_aelse_acc_nl;
  wire Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_nl;
  wire[9:0] operator_9_false_1_acc_nl;
  wire[10:0] nl_operator_9_false_1_acc_nl;
  wire[8:0] operator_9_false_acc_nl;
  wire[9:0] nl_operator_9_false_acc_nl;
  wire[8:0] Tensor_weight_y_COLUMN_if_4_mux_1_nl;
  wire[8:0] Tensor_weight_y_ROW_acc_nl;
  wire[9:0] nl_Tensor_weight_y_ROW_acc_nl;
  wire Tensor_weight_y_ROW_not_17_nl;
  wire[10:0] Tensor_weight_y_COLUMN_if_4_mux_nl;
  wire Tensor_weight_y_ROW_Tensor_weight_y_ROW_Tensor_weight_y_ROW_Tensor_weight_y_ROW_not_nl;
  wire[9:0] operator_9_false_acc_nl_1;
  wire[10:0] nl_operator_9_false_acc_nl_1;
  wire[94:0] Tensor_weight_y_COLUMN_if_3_acc_39_nl;
  wire[96:0] nl_Tensor_weight_y_COLUMN_if_3_acc_39_nl;
  wire[63:0] Tensor_weight_y_COLUMN_if_3_acc_37_nl;
  wire[64:0] nl_Tensor_weight_y_COLUMN_if_3_acc_37_nl;
  wire[383:0] out_product0_val_mux_nl;
  wire and_120_nl;
  wire[94:0] Tensor_weight_y_COLUMN_if_3_acc_nl;
  wire[95:0] nl_Tensor_weight_y_COLUMN_if_3_acc_nl;
  wire[93:0] Tensor_weight_y_COLUMN_if_3_acc_50_nl;
  wire[94:0] nl_Tensor_weight_y_COLUMN_if_3_acc_50_nl;
  wire[63:0] Tensor_weight_y_COLUMN_if_3_mux_18_nl;
  wire[29:0] Tensor_weight_y_COLUMN_if_3_mux_19_nl;
  wire[94:0] Tensor_weight_y_COLUMN_if_3_acc_52_nl;
  wire[95:0] nl_Tensor_weight_y_COLUMN_if_3_acc_52_nl;
  wire[93:0] Tensor_weight_y_COLUMN_if_3_acc_51_nl;
  wire[94:0] nl_Tensor_weight_y_COLUMN_if_3_acc_51_nl;
  wire[63:0] Tensor_weight_y_COLUMN_if_3_mux_20_nl;
  wire[29:0] Tensor_weight_y_COLUMN_if_3_mux_21_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [383:0] nl_OpticalFlow_tensor_weight_y_run_tensor_y_rsci_inst_tensor_y_rsci_idat;
  assign nl_OpticalFlow_tensor_weight_y_run_tensor_y_rsci_inst_tensor_y_rsci_idat
      = {tensor_y_rsci_idat_383_320 , tensor_y_rsci_idat_319_256 , tensor_y_rsci_idat_255_192
      , tensor_y_rsci_idat_191_128 , tensor_y_rsci_idat_127_64 , tensor_y_rsci_idat_63_0};
  OpticalFlow_tensor_weight_y_run_out_product_rsci OpticalFlow_tensor_weight_y_run_out_product_rsci_inst
      (
      .out_product_rsc_dat(out_product_rsc_dat),
      .out_product_rsc_vld(out_product_rsc_vld),
      .out_product_rsc_rdy(out_product_rsc_rdy),
      .run_wen(run_wen),
      .out_product_rsci_oswt(reg_out_product_rsci_iswt0_cse),
      .out_product_rsci_wen_comp(out_product_rsci_wen_comp),
      .out_product_rsci_idat_mxwt(out_product_rsci_idat_mxwt)
    );
  OpticalFlow_tensor_weight_y_run_tensor_y_rsci OpticalFlow_tensor_weight_y_run_tensor_y_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_y_rsc_dat(tensor_y_rsc_dat),
      .tensor_y_rsc_vld(tensor_y_rsc_vld),
      .tensor_y_rsc_rdy(tensor_y_rsc_rdy),
      .run_wen(run_wen),
      .tensor_y_rsci_oswt(reg_tensor_y_rsci_iswt0_cse),
      .tensor_y_rsci_wen_comp(tensor_y_rsci_wen_comp),
      .tensor_y_rsci_idat(nl_OpticalFlow_tensor_weight_y_run_tensor_y_rsci_inst_tensor_y_rsci_idat[383:0])
    );
  OpticalFlow_tensor_weight_y_run_wait_dp OpticalFlow_tensor_weight_y_run_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z),
      .run_wen(run_wen),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg)
    );
  OpticalFlow_tensor_weight_y_run_staller OpticalFlow_tensor_weight_y_run_staller_inst
      (
      .run_wen(run_wen),
      .out_product_rsci_wen_comp(out_product_rsci_wen_comp),
      .tensor_y_rsci_wen_comp(tensor_y_rsci_wen_comp)
    );
  OpticalFlow_tensor_weight_y_run_run_fsm OpticalFlow_tensor_weight_y_run_run_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign line_buf1_rsci_clken_d = run_wen;
  assign Tensor_weight_y_COLUMN_if_3_or_itm = and_40_cse | (main_stage_0_3 & Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_and_itm_1
      & (fsm_output[2]));
  assign Tensor_weight_y_COLUMN_if_3_and_cse = run_wen & Tensor_weight_y_COLUMN_if_3_or_itm;
  assign Tensor_weight_y_COLUMN_if_3_and_6_cse = run_wen & (fsm_output[2]);
  assign rdbuf0_and_cse = run_wen & (~ (Tensor_weight_y_COLUMN_x_lpi_1_dfm[0])) &
      (fsm_output[2]);
  assign Tensor_weight_y_COLUMN_qelse_1_and_cse = run_wen & (Tensor_weight_y_COLUMN_x_lpi_1_dfm_1_0
      | (fsm_output[2]));
  assign and_37_cse = Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1
      & Tensor_weight_y_ROW_equal_1_tmp;
  assign out_product0_val_lpi_1_dfm_mx1 = MUX_v_384_2_2(out_product_rsci_idat_mxwt,
      out_product0_val_lpi_1, Tensor_weight_y_COLUMN_if_slc_Tensor_weight_y_COLUMN_acc_9_svs);
  assign exitL_exit_Tensor_weight_y_ROW_sva_mx0 = and_37_cse | (~ main_stage_0_2);
  assign Tensor_weight_y_ROW_equal_1_tmp = Tensor_weight_y_ROW_y_lpi_1_dfm == heightIn;
  assign Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_mx1_383_192 = MUX_v_192_2_2(Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_383_192,
      (rdbuf0_lpi_1[767:576]), Tensor_weight_y_COLUMN_x_lpi_1_dfm_1_0);
  assign Tensor_weight_y_COLUMN_qr_lpi_1_dfm_mx1_383_192 = MUX_v_192_2_2(Tensor_weight_y_COLUMN_qr_lpi_1_dfm_383_192,
      (rdbuf1_lpi_1_767_384[383:192]), Tensor_weight_y_COLUMN_x_lpi_1_dfm_1_0);
  assign nl_Tensor_weight_y_ROW_acc_nl = Tensor_weight_y_ROW_y_lpi_1_dfm + 9'b000000001;
  assign Tensor_weight_y_ROW_acc_nl = nl_Tensor_weight_y_ROW_acc_nl[8:0];
  assign Tensor_weight_y_COLUMN_if_4_mux_1_nl = MUX_v_9_2_2(Tensor_weight_y_ROW_y_lpi_1_dfm,
      Tensor_weight_y_ROW_acc_nl, Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1);
  assign Tensor_weight_y_ROW_not_17_nl = ~ exitL_exit_Tensor_weight_y_ROW_sva_mx0;
  assign Tensor_weight_y_ROW_y_lpi_1_dfm_mx0w0 = MUX_v_9_2_2(9'b000000000, Tensor_weight_y_COLUMN_if_4_mux_1_nl,
      Tensor_weight_y_ROW_not_17_nl);
  assign Tensor_weight_y_COLUMN_if_4_mux_nl = MUX_v_11_2_2(Tensor_weight_y_COLUMN_x_sva_2_1,
      ({{10{Tensor_weight_y_ROW_equal_1_tmp}}, Tensor_weight_y_ROW_equal_1_tmp}),
      Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1);
  assign Tensor_weight_y_ROW_Tensor_weight_y_ROW_Tensor_weight_y_ROW_Tensor_weight_y_ROW_not_nl
      = ~ exitL_exit_Tensor_weight_y_ROW_sva_mx0;
  assign Tensor_weight_y_COLUMN_x_lpi_1_dfm_2 = MUX_v_11_2_2(11'b00000000000, Tensor_weight_y_COLUMN_if_4_mux_nl,
      Tensor_weight_y_ROW_Tensor_weight_y_ROW_Tensor_weight_y_ROW_Tensor_weight_y_ROW_not_nl);
  assign nl_operator_9_false_acc_nl_1 = ({1'b1 , heightIn}) + conv_u2s_9_10(~ Tensor_weight_y_ROW_y_lpi_1_dfm_mx0w0);
  assign operator_9_false_acc_nl_1 = nl_operator_9_false_acc_nl_1[9:0];
  assign operator_9_false_acc_itm_9_1 = readslicef_10_1_9(operator_9_false_acc_nl_1);
  assign nl_operator_11_false_acc_psp_sva_1 = conv_u2s_11_12(widthIn) + 12'b111111111111;
  assign operator_11_false_acc_psp_sva_1 = nl_operator_11_false_acc_psp_sva_1[11:0];
  assign nl_Tensor_weight_y_COLUMN_if_3_acc_37_nl = (Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg[93:30])
      + 64'b0000000000000000000000000000000000000000000000000000000000000001;
  assign Tensor_weight_y_COLUMN_if_3_acc_37_nl = nl_Tensor_weight_y_COLUMN_if_3_acc_37_nl[63:0];
  assign nl_Tensor_weight_y_COLUMN_if_3_acc_39_nl = conv_s2s_94_95({Tensor_weight_y_COLUMN_if_3_acc_37_nl
      , (Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z_oreg[29:0])}) + conv_s2s_94_95(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z_oreg)
      + conv_s2s_94_95({Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z_oreg , 1'b0});
  assign Tensor_weight_y_COLUMN_if_3_acc_39_nl = nl_Tensor_weight_y_COLUMN_if_3_acc_39_nl[94:0];
  assign Tensor_weight_y_COLUMN_if_3_acc_39_itm_94_31_1 = readslicef_95_64_31(Tensor_weight_y_COLUMN_if_3_acc_39_nl);
  assign nl_Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_9_93_30
      = (Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg[93:30]) + 64'b0000000000000000000000000000000000000000000000000000000000000001;
  assign Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_9_93_30 = nl_Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_9_93_30[63:0];
  assign nl_Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_11_93_30
      = (Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg[93:30]) + 64'b0000000000000000000000000000000000000000000000000000000000000001;
  assign Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_11_93_30 =
      nl_Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_11_93_30[63:0];
  assign Tensor_weight_y_COLUMN_if_4_mux_1_tmp_0 = MUX_s_1_2_2((Tensor_weight_y_COLUMN_x_sva_2_1[0]),
      Tensor_weight_y_ROW_equal_1_tmp, Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1);
  assign and_40_cse = main_stage_0_3 & (~ Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_and_itm_1)
      & (~ operator_9_false_1_slc_operator_9_false_1_acc_9_itm) & (fsm_output[1]);
  assign line_buf1_rsci_adr_d = Tensor_weight_y_COLUMN_x_lpi_1_dfm_2[9:1];
  assign line_buf1_rsci_d_d = rdbuf0_lpi_1;
  assign line_buf1_rsci_we_d_pff = (~(Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1
      & Tensor_weight_y_ROW_equal_1_tmp)) & main_stage_0_2 & Tensor_weight_y_COLUMN_if_4_mux_1_tmp_0
      & (fsm_output[1]);
  assign line_buf1_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff = (and_37_cse | (~(main_stage_0_2
      & Tensor_weight_y_COLUMN_if_4_mux_1_tmp_0))) & (fsm_output[1]);
  assign line_buf0_rsci_adr_d = MUX_v_9_2_2((Tensor_weight_y_COLUMN_x_lpi_1_dfm_2[9:1]),
      (Tensor_weight_y_COLUMN_x_lpi_1_dfm[9:1]), fsm_output[2]);
  assign and_120_nl = (~ Tensor_weight_y_COLUMN_if_slc_Tensor_weight_y_COLUMN_acc_9_svs)
      & (fsm_output[2]);
  assign out_product0_val_mux_nl = MUX_v_384_2_2(out_product0_val_lpi_1, out_product_rsci_idat_mxwt,
      and_120_nl);
  assign line_buf0_rsci_d_d = {out_product0_val_mux_nl , wrbuf0_383_320_lpi_1_dfm_2
      , wrbuf0_319_256_lpi_1_dfm_2 , wrbuf0_255_192_lpi_1_dfm_2 , wrbuf0_191_128_lpi_1_dfm_2
      , wrbuf0_127_64_lpi_1_dfm_2 , wrbuf0_63_0_lpi_1_dfm_2};
  assign line_buf0_rsci_we_d_pff = (Tensor_weight_y_COLUMN_x_lpi_1_dfm[0]) & (fsm_output[2]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      tensor_y_rsci_idat_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_127_64 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_191_128 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_255_192 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_319_256 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_383_320 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      tensor_y_rsci_idat_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_127_64 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_191_128 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_255_192 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_319_256 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tensor_y_rsci_idat_383_320 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( Tensor_weight_y_COLUMN_if_3_and_cse ) begin
      tensor_y_rsci_idat_63_0 <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          Tensor_weight_y_COLUMN_if_3_acc_39_itm_94_31_1, Tensor_weight_y_COLUMN_if_3_not_6_nl);
      tensor_y_rsci_idat_127_64 <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          z_out_94_31, Tensor_weight_y_COLUMN_if_3_not_7_nl);
      tensor_y_rsci_idat_191_128 <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          z_out_1_94_31, Tensor_weight_y_COLUMN_if_3_not_8_nl);
      tensor_y_rsci_idat_255_192 <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          Tensor_weight_y_COLUMN_if_3_slc_94_31_3_itm, Tensor_weight_y_COLUMN_if_3_not_9_nl);
      tensor_y_rsci_idat_319_256 <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          Tensor_weight_y_COLUMN_if_3_slc_94_31_4_itm, Tensor_weight_y_COLUMN_if_3_not_10_nl);
      tensor_y_rsci_idat_383_320 <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          Tensor_weight_y_COLUMN_if_3_slc_94_31_5_itm, Tensor_weight_y_COLUMN_if_3_not_11_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_tensor_y_rsci_iswt0_cse <= 1'b0;
      reg_out_product_rsci_iswt0_cse <= 1'b0;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      out_product0_val_lpi_1 <= 384'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_x_lpi_1_dfm_1_0 <= 1'b0;
      Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1
          <= 1'b0;
      Tensor_weight_y_COLUMN_x_sva_2_1 <= 11'b00000000000;
      operator_9_false_slc_operator_9_false_acc_8_svs_1 <= 1'b0;
      Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_383_192 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_qr_lpi_1_dfm_383_192 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_slc_94_31_3_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_slc_94_31_4_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_slc_94_31_5_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_x_lpi_1_dfm <= 11'b00000000000;
      Tensor_weight_y_COLUMN_if_slc_Tensor_weight_y_COLUMN_acc_9_svs <= 1'b0;
      operator_9_false_slc_operator_9_false_acc_8_svs <= 1'b0;
    end
    else if ( rst ) begin
      reg_tensor_y_rsci_iswt0_cse <= 1'b0;
      reg_out_product_rsci_iswt0_cse <= 1'b0;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      out_product0_val_lpi_1 <= 384'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_x_lpi_1_dfm_1_0 <= 1'b0;
      Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1
          <= 1'b0;
      Tensor_weight_y_COLUMN_x_sva_2_1 <= 11'b00000000000;
      operator_9_false_slc_operator_9_false_acc_8_svs_1 <= 1'b0;
      Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_383_192 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_qr_lpi_1_dfm_383_192 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_slc_94_31_3_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_slc_94_31_4_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_if_3_slc_94_31_5_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_x_lpi_1_dfm <= 11'b00000000000;
      Tensor_weight_y_COLUMN_if_slc_Tensor_weight_y_COLUMN_acc_9_svs <= 1'b0;
      operator_9_false_slc_operator_9_false_acc_8_svs <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_tensor_y_rsci_iswt0_cse <= Tensor_weight_y_COLUMN_if_3_or_itm;
      reg_out_product_rsci_iswt0_cse <= (~ operator_9_false_acc_itm_9_1) & (fsm_output[1]);
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b <= MUX_v_64_2_2((Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_mx1_383_192[191:128]),
          (Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_191_0[191:128]), fsm_output[2]);
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b <= MUX_v_64_2_2((Tensor_weight_y_COLUMN_qr_lpi_1_dfm_mx1_383_192[191:128]),
          (Tensor_weight_y_COLUMN_qr_lpi_1_dfm_191_0[127:64]), fsm_output[2]);
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b <= MUX_v_64_2_2((out_product0_val_lpi_1_dfm_1[319:256]),
          (out_product0_val_lpi_1_dfm_1[127:64]), fsm_output[2]);
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b <= MUX_v_64_2_2((Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_mx1_383_192[127:64]),
          (Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_191_0[127:64]), fsm_output[2]);
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b <= MUX_v_64_2_2((Tensor_weight_y_COLUMN_qr_lpi_1_dfm_mx1_383_192[127:64]),
          (Tensor_weight_y_COLUMN_qr_lpi_1_dfm_191_0[191:128]), fsm_output[2]);
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b <= MUX_v_64_2_2((out_product0_val_lpi_1_dfm_1[255:192]),
          (out_product0_val_lpi_1_dfm_1[63:0]), fsm_output[2]);
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b <= MUX_v_64_2_2((Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_mx1_383_192[63:0]),
          (Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_191_0[63:0]), fsm_output[2]);
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b <= MUX_v_64_2_2((Tensor_weight_y_COLUMN_qr_lpi_1_dfm_mx1_383_192[63:0]),
          (Tensor_weight_y_COLUMN_qr_lpi_1_dfm_191_0[63:0]), fsm_output[2]);
      Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b <= MUX_v_64_2_2((out_product0_val_lpi_1_dfm_1[383:320]),
          (out_product0_val_lpi_1_dfm_1[191:128]), fsm_output[2]);
      out_product0_val_lpi_1 <= out_product0_val_lpi_1_dfm_1;
      Tensor_weight_y_COLUMN_x_lpi_1_dfm_1_0 <= Tensor_weight_y_COLUMN_x_lpi_1_dfm[0];
      Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1
          <= MUX_s_1_2_2(Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_and_nl,
          Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_nl,
          fsm_output[2]);
      Tensor_weight_y_COLUMN_x_sva_2_1 <= nl_Tensor_weight_y_COLUMN_x_sva_2_1[10:0];
      operator_9_false_slc_operator_9_false_acc_8_svs_1 <= operator_9_false_slc_operator_9_false_acc_8_svs;
      Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_383_192 <= line_buf0_rsci_q_d[383:192];
      Tensor_weight_y_COLUMN_qr_lpi_1_dfm_383_192 <= line_buf1_rsci_q_d[383:192];
      Tensor_weight_y_COLUMN_if_3_slc_94_31_3_itm <= Tensor_weight_y_COLUMN_if_3_acc_39_itm_94_31_1;
      Tensor_weight_y_COLUMN_if_3_slc_94_31_4_itm <= z_out_94_31;
      Tensor_weight_y_COLUMN_if_3_slc_94_31_5_itm <= z_out_1_94_31;
      Tensor_weight_y_COLUMN_x_lpi_1_dfm <= Tensor_weight_y_COLUMN_x_lpi_1_dfm_2;
      Tensor_weight_y_COLUMN_if_slc_Tensor_weight_y_COLUMN_acc_9_svs <= operator_9_false_acc_itm_9_1;
      operator_9_false_slc_operator_9_false_acc_8_svs <= readslicef_9_1_8(operator_9_false_acc_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_and_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
    end
    else if ( rst ) begin
      Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_and_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
    end
    else if ( Tensor_weight_y_COLUMN_if_3_and_6_cse ) begin
      Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_and_itm_1 <= Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_svs_1;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      out_product0_val_lpi_1_dfm_1 <= 384'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      out_product0_val_lpi_1_dfm_1 <= 384'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~ (fsm_output[1])) ) begin
      out_product0_val_lpi_1_dfm_1 <= MUX_v_384_2_2(out_product_rsci_idat_mxwt, out_product0_val_lpi_1,
          and_122_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rdbuf0_lpi_1 <= 768'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_383_320_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_319_256_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_255_192_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_191_128_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_127_64_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_63_0_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf1_lpi_1_767_384 <= 384'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      rdbuf0_lpi_1 <= 768'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_383_320_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_319_256_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_255_192_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_191_128_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_127_64_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      wrbuf0_63_0_lpi_1_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf1_lpi_1_767_384 <= 384'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rdbuf0_and_cse ) begin
      rdbuf0_lpi_1 <= line_buf0_rsci_q_d;
      wrbuf0_383_320_lpi_1_dfm_2 <= out_product0_val_lpi_1_dfm_mx1[383:320];
      wrbuf0_319_256_lpi_1_dfm_2 <= out_product0_val_lpi_1_dfm_mx1[319:256];
      wrbuf0_255_192_lpi_1_dfm_2 <= out_product0_val_lpi_1_dfm_mx1[255:192];
      wrbuf0_191_128_lpi_1_dfm_2 <= out_product0_val_lpi_1_dfm_mx1[191:128];
      wrbuf0_127_64_lpi_1_dfm_2 <= out_product0_val_lpi_1_dfm_mx1[127:64];
      wrbuf0_63_0_lpi_1_dfm_2 <= out_product0_val_lpi_1_dfm_mx1[63:0];
      rdbuf1_lpi_1_767_384 <= line_buf1_rsci_q_d[767:384];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_191_0 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_qr_lpi_1_dfm_191_0 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_191_0 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      Tensor_weight_y_COLUMN_qr_lpi_1_dfm_191_0 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( Tensor_weight_y_COLUMN_qelse_1_and_cse ) begin
      Tensor_weight_y_COLUMN_qr_1_lpi_1_dfm_191_0 <= MUX_v_192_2_2((rdbuf0_lpi_1[575:384]),
          (line_buf0_rsci_q_d[191:0]), fsm_output[2]);
      Tensor_weight_y_COLUMN_qr_lpi_1_dfm_191_0 <= MUX_v_192_2_2((rdbuf1_lpi_1_767_384[191:0]),
          (line_buf1_rsci_q_d[191:0]), fsm_output[2]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      Tensor_weight_y_ROW_y_lpi_1_dfm <= 9'b000000000;
    end
    else if ( rst ) begin
      Tensor_weight_y_ROW_y_lpi_1_dfm <= 9'b000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      Tensor_weight_y_ROW_y_lpi_1_dfm <= Tensor_weight_y_ROW_y_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm <= 1'b0;
    end
    else if ( rst ) begin
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm <= 1'b0;
    end
    else if ( run_wen & (~ (fsm_output[2])) ) begin
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm <= readslicef_10_1_9(operator_9_false_1_acc_nl);
    end
  end
  assign Tensor_weight_y_COLUMN_if_3_not_6_nl = ~ and_40_cse;
  assign Tensor_weight_y_COLUMN_if_3_not_7_nl = ~ and_40_cse;
  assign Tensor_weight_y_COLUMN_if_3_not_8_nl = ~ and_40_cse;
  assign Tensor_weight_y_COLUMN_if_3_not_9_nl = ~ and_40_cse;
  assign Tensor_weight_y_COLUMN_if_3_not_10_nl = ~ and_40_cse;
  assign Tensor_weight_y_COLUMN_if_3_not_11_nl = ~ and_40_cse;
  assign nl_Tensor_weight_y_COLUMN_aelse_acc_nl = ({1'b1 , Tensor_weight_y_ROW_y_lpi_1_dfm})
      + conv_u2u_9_10(~ heightIn) + 10'b0000000001;
  assign Tensor_weight_y_COLUMN_aelse_acc_nl = nl_Tensor_weight_y_COLUMN_aelse_acc_nl[9:0];
  assign Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_and_nl = (readslicef_10_1_9(Tensor_weight_y_COLUMN_aelse_acc_nl))
      & (~ operator_9_false_slc_operator_9_false_acc_8_svs_1);
  assign Tensor_weight_y_COLUMN_Tensor_weight_y_COLUMN_if_4_Tensor_weight_y_COLUMN_if_4_nor_nl
      = ~((Tensor_weight_y_COLUMN_x_lpi_1_dfm != (operator_11_false_acc_psp_sva_1[10:0]))
      | (operator_11_false_acc_psp_sva_1[11]));
  assign nl_Tensor_weight_y_COLUMN_x_sva_2_1  = Tensor_weight_y_COLUMN_x_lpi_1_dfm
      + 11'b00000000001;
  assign nl_operator_9_false_acc_nl = conv_u2u_8_9(Tensor_weight_y_ROW_y_lpi_1_dfm_mx0w0[8:1])
      + 9'b111111111;
  assign operator_9_false_acc_nl = nl_operator_9_false_acc_nl[8:0];
  assign and_122_nl = Tensor_weight_y_COLUMN_if_slc_Tensor_weight_y_COLUMN_acc_9_svs
      & (fsm_output[2]);
  assign nl_operator_9_false_1_acc_nl = conv_u2s_9_10(Tensor_weight_y_ROW_y_lpi_1_dfm)
      + 10'b1111111111;
  assign operator_9_false_1_acc_nl = nl_operator_9_false_1_acc_nl[9:0];
  assign nl_Tensor_weight_y_COLUMN_if_3_acc_50_nl = conv_s2s_93_94(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg[93:1])
      + conv_s2s_93_94(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z_oreg);
  assign Tensor_weight_y_COLUMN_if_3_acc_50_nl = nl_Tensor_weight_y_COLUMN_if_3_acc_50_nl[93:0];
  assign Tensor_weight_y_COLUMN_if_3_mux_18_nl = MUX_v_64_2_2(Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_9_93_30,
      Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_11_93_30, fsm_output[1]);
  assign Tensor_weight_y_COLUMN_if_3_mux_19_nl = MUX_v_30_2_2((Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg[29:0]),
      (Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg[29:0]), fsm_output[1]);
  assign nl_Tensor_weight_y_COLUMN_if_3_acc_nl = ({Tensor_weight_y_COLUMN_if_3_acc_50_nl
      , (Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z_oreg[0])}) + conv_s2u_94_95({Tensor_weight_y_COLUMN_if_3_mux_18_nl
      , Tensor_weight_y_COLUMN_if_3_mux_19_nl});
  assign Tensor_weight_y_COLUMN_if_3_acc_nl = nl_Tensor_weight_y_COLUMN_if_3_acc_nl[94:0];
  assign z_out_94_31 = readslicef_95_64_31(Tensor_weight_y_COLUMN_if_3_acc_nl);
  assign nl_Tensor_weight_y_COLUMN_if_3_acc_51_nl = conv_s2s_93_94(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg[93:1])
      + conv_s2s_93_94(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z_oreg);
  assign Tensor_weight_y_COLUMN_if_3_acc_51_nl = nl_Tensor_weight_y_COLUMN_if_3_acc_51_nl[93:0];
  assign Tensor_weight_y_COLUMN_if_3_mux_20_nl = MUX_v_64_2_2(Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_11_93_30,
      Tensor_weight_y_COLUMN_if_3_Tensor_weight_y_COLUMN_if_3_conc_9_93_30, fsm_output[1]);
  assign Tensor_weight_y_COLUMN_if_3_mux_21_nl = MUX_v_30_2_2((Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z_oreg[29:0]),
      (Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z_oreg[29:0]), fsm_output[1]);
  assign nl_Tensor_weight_y_COLUMN_if_3_acc_52_nl = ({Tensor_weight_y_COLUMN_if_3_acc_51_nl
      , (Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z_oreg[0])}) + conv_s2u_94_95({Tensor_weight_y_COLUMN_if_3_mux_20_nl
      , Tensor_weight_y_COLUMN_if_3_mux_21_nl});
  assign Tensor_weight_y_COLUMN_if_3_acc_52_nl = nl_Tensor_weight_y_COLUMN_if_3_acc_52_nl[94:0];
  assign z_out_1_94_31 = readslicef_95_64_31(Tensor_weight_y_COLUMN_if_3_acc_52_nl);

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [191:0] MUX_v_192_2_2;
    input [191:0] input_0;
    input [191:0] input_1;
    input  sel;
    reg [191:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_192_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input  sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [383:0] MUX_v_384_2_2;
    input [383:0] input_0;
    input [383:0] input_1;
    input  sel;
    reg [383:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_384_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [63:0] readslicef_95_64_31;
    input [94:0] vector;
    reg [94:0] tmp;
  begin
    tmp = vector >> 31;
    readslicef_95_64_31 = tmp[63:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [93:0] conv_s2s_93_94 ;
    input [92:0]  vector ;
  begin
    conv_s2s_93_94 = {vector[92], vector};
  end
  endfunction


  function automatic [94:0] conv_s2s_94_95 ;
    input [93:0]  vector ;
  begin
    conv_s2s_94_95 = {vector[93], vector};
  end
  endfunction


  function automatic [94:0] conv_s2u_94_95 ;
    input [93:0]  vector ;
  begin
    conv_s2u_94_95 = {vector[93], vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y_struct
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y_struct (
  clk, rst, arst_n, out_product_rsc_dat_val, out_product_rsc_vld, out_product_rsc_rdy,
      tensor_y_rsc_dat_val, tensor_y_rsc_vld, tensor_y_rsc_rdy, widthIn, heightIn,
      line_buf1_rsc_clken, line_buf1_rsc_q, line_buf1_rsc_we, line_buf1_rsc_d, line_buf1_rsc_adr,
      line_buf0_rsc_clken, line_buf0_rsc_q, line_buf0_rsc_we, line_buf0_rsc_d, line_buf0_rsc_adr
);
  input clk;
  input rst;
  input arst_n;
  input [383:0] out_product_rsc_dat_val;
  input out_product_rsc_vld;
  output out_product_rsc_rdy;
  output [383:0] tensor_y_rsc_dat_val;
  output tensor_y_rsc_vld;
  input tensor_y_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  output line_buf1_rsc_clken;
  input [767:0] line_buf1_rsc_q;
  output line_buf1_rsc_we;
  output [767:0] line_buf1_rsc_d;
  output [8:0] line_buf1_rsc_adr;
  output line_buf0_rsc_clken;
  input [767:0] line_buf0_rsc_q;
  output line_buf0_rsc_we;
  output [767:0] line_buf0_rsc_d;
  output [8:0] line_buf0_rsc_adr;


  // Interconnect Declarations
  wire [8:0] line_buf1_rsci_adr_d;
  wire line_buf1_rsci_clken_d;
  wire [767:0] line_buf1_rsci_d_d;
  wire [767:0] line_buf1_rsci_q_d;
  wire [8:0] line_buf0_rsci_adr_d;
  wire [767:0] line_buf0_rsci_d_d;
  wire [767:0] line_buf0_rsci_q_d;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b;
  wire [63:0] Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b;
  wire [383:0] tensor_y_rsc_dat;
  wire line_buf1_rsci_we_d_iff;
  wire line_buf1_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff;
  wire line_buf0_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [94:0] nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z;
  assign nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b);
  wire [94:0] nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z;
  assign nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b);
  wire[92:0] mul_2_nl;
  wire signed [93:0] nl_mul_2_nl;
  wire [93:0] nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z;
  assign nl_mul_2_nl = $signed(30'b010110011110111011001011111111) * $signed(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b);
  assign mul_2_nl = nl_mul_2_nl[92:0];
  assign nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z
      = signext_94_93(mul_2_nl);
  wire [94:0] nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z;
  assign nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b);
  wire [94:0] nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z;
  assign nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b);
  wire[92:0] mul_5_nl;
  wire signed [93:0] nl_mul_5_nl;
  wire [93:0] nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z;
  assign nl_mul_5_nl = $signed(30'b010110011110111011001011111111) * $signed(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b);
  assign mul_5_nl = nl_mul_5_nl[92:0];
  assign nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z
      = signext_94_93(mul_5_nl);
  wire [94:0] nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z;
  assign nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b);
  wire [94:0] nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z;
  assign nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z
      = $signed(31'b0101001100000101010100110010011) * $signed(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b);
  wire[92:0] mul_8_nl;
  wire signed [93:0] nl_mul_8_nl;
  wire [93:0] nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z;
  assign nl_mul_8_nl = $signed(30'b010110011110111011001011111111) * $signed(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b);
  assign mul_8_nl = nl_mul_8_nl[92:0];
  assign nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z
      = signext_94_93(mul_8_nl);
  OpticalFlow_tensor_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_5_9_768_512_1_512_768_1_gen
      line_buf1_rsci (
      .clken(line_buf1_rsc_clken),
      .q(line_buf1_rsc_q),
      .we(line_buf1_rsc_we),
      .d(line_buf1_rsc_d),
      .adr(line_buf1_rsc_adr),
      .adr_d(line_buf1_rsci_adr_d),
      .clken_d(line_buf1_rsci_clken_d),
      .d_d(line_buf1_rsci_d_d),
      .q_d(line_buf1_rsci_q_d),
      .we_d(line_buf1_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf1_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf1_rsci_we_d_iff)
    );
  OpticalFlow_tensor_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_6_9_768_512_1_512_768_1_gen
      line_buf0_rsci (
      .clken(line_buf0_rsc_clken),
      .q(line_buf0_rsc_q),
      .we(line_buf0_rsc_we),
      .d(line_buf0_rsc_d),
      .adr(line_buf0_rsc_adr),
      .adr_d(line_buf0_rsci_adr_d),
      .clken_d(line_buf1_rsci_clken_d),
      .d_d(line_buf0_rsci_d_d),
      .q_d(line_buf0_rsci_q_d),
      .we_d(line_buf0_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf1_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf0_rsci_we_d_iff)
    );
  OpticalFlow_tensor_weight_y_run OpticalFlow_tensor_weight_y_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .out_product_rsc_dat(out_product_rsc_dat_val),
      .out_product_rsc_vld(out_product_rsc_vld),
      .out_product_rsc_rdy(out_product_rsc_rdy),
      .tensor_y_rsc_dat(tensor_y_rsc_dat),
      .tensor_y_rsc_vld(tensor_y_rsc_vld),
      .tensor_y_rsc_rdy(tensor_y_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .line_buf1_rsci_adr_d(line_buf1_rsci_adr_d),
      .line_buf1_rsci_clken_d(line_buf1_rsci_clken_d),
      .line_buf1_rsci_d_d(line_buf1_rsci_d_d),
      .line_buf1_rsci_q_d(line_buf1_rsci_q_d),
      .line_buf0_rsci_adr_d(line_buf0_rsci_adr_d),
      .line_buf0_rsci_d_d(line_buf0_rsci_d_d),
      .line_buf0_rsci_q_d(line_buf0_rsci_q_d),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_b),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z(nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_z[93:0]),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_b),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z(nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_1_z[93:0]),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_b),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z(nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_2_z[93:0]),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_b),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z(nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_3_z[93:0]),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_b),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z(nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_4_z[93:0]),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_b),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z(nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_5_z[93:0]),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_b),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z(nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_6_z[93:0]),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_b),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z(nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_7_z[93:0]),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b(Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_b),
      .Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z(nl_OpticalFlow_tensor_weight_y_run_inst_Tensor_weight_y_COLUMN_if_3_mul_15_cmp_8_z[93:0]),
      .line_buf1_rsci_we_d_pff(line_buf1_rsci_we_d_iff),
      .line_buf1_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff(line_buf1_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .line_buf0_rsci_we_d_pff(line_buf0_rsci_we_d_iff)
    );
  assign tensor_y_rsc_dat_val = tensor_y_rsc_dat;

  function automatic [93:0] signext_94_93;
    input [92:0] vector;
  begin
    signext_94_93= {{1{vector[92]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_tensor_weight_y
// ------------------------------------------------------------------


module OpticalFlow_tensor_weight_y (
  clk, rst, arst_n, out_product_rsc_dat, out_product_rsc_vld, out_product_rsc_rdy,
      tensor_y_rsc_dat, tensor_y_rsc_vld, tensor_y_rsc_rdy, widthIn, heightIn, line_buf1_rsc_clken,
      line_buf1_rsc_q, line_buf1_rsc_we, line_buf1_rsc_d, line_buf1_rsc_adr, line_buf0_rsc_clken,
      line_buf0_rsc_q, line_buf0_rsc_we, line_buf0_rsc_d, line_buf0_rsc_adr
);
  input clk;
  input rst;
  input arst_n;
  input [383:0] out_product_rsc_dat;
  input out_product_rsc_vld;
  output out_product_rsc_rdy;
  output [383:0] tensor_y_rsc_dat;
  output tensor_y_rsc_vld;
  input tensor_y_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  output line_buf1_rsc_clken;
  input [767:0] line_buf1_rsc_q;
  output line_buf1_rsc_we;
  output [767:0] line_buf1_rsc_d;
  output [8:0] line_buf1_rsc_adr;
  output line_buf0_rsc_clken;
  input [767:0] line_buf0_rsc_q;
  output line_buf0_rsc_we;
  output [767:0] line_buf0_rsc_d;
  output [8:0] line_buf0_rsc_adr;


  // Interconnect Declarations
  wire [383:0] tensor_y_rsc_dat_val;


  // Interconnect Declarations for Component Instantiations 
  OpticalFlow_tensor_weight_y_struct OpticalFlow_tensor_weight_y_struct_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .out_product_rsc_dat_val(out_product_rsc_dat),
      .out_product_rsc_vld(out_product_rsc_vld),
      .out_product_rsc_rdy(out_product_rsc_rdy),
      .tensor_y_rsc_dat_val(tensor_y_rsc_dat_val),
      .tensor_y_rsc_vld(tensor_y_rsc_vld),
      .tensor_y_rsc_rdy(tensor_y_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .line_buf1_rsc_clken(line_buf1_rsc_clken),
      .line_buf1_rsc_q(line_buf1_rsc_q),
      .line_buf1_rsc_we(line_buf1_rsc_we),
      .line_buf1_rsc_d(line_buf1_rsc_d),
      .line_buf1_rsc_adr(line_buf1_rsc_adr),
      .line_buf0_rsc_clken(line_buf0_rsc_clken),
      .line_buf0_rsc_q(line_buf0_rsc_q),
      .line_buf0_rsc_we(line_buf0_rsc_we),
      .line_buf0_rsc_d(line_buf0_rsc_d),
      .line_buf0_rsc_adr(line_buf0_rsc_adr)
    );
  assign tensor_y_rsc_dat = tensor_y_rsc_dat_val;
endmodule




//------> ../OpticalFlow_outer_product.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Sun Jun 16 21:08:19 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module OpticalFlow_outer_product_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for OpticalFlow_outer_product_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : OpticalFlow_outer_product_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product_run_staller
// ------------------------------------------------------------------


module OpticalFlow_outer_product_run_staller (
  run_wen, filtered_gradient_rsci_wen_comp, out_product_rsci_wen_comp
);
  output run_wen;
  input filtered_gradient_rsci_wen_comp;
  input out_product_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = filtered_gradient_rsci_wen_comp & out_product_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product_run_out_product_rsci_out_product_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_outer_product_run_out_product_rsci_out_product_wait_dp (
  clk, rst, arst_n, out_product_rsci_oswt, out_product_rsci_wen_comp, out_product_rsci_biwt,
      out_product_rsci_bdwt, out_product_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input out_product_rsci_oswt;
  output out_product_rsci_wen_comp;
  input out_product_rsci_biwt;
  input out_product_rsci_bdwt;
  output out_product_rsci_bcwt;
  reg out_product_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign out_product_rsci_wen_comp = (~ out_product_rsci_oswt) | out_product_rsci_biwt
      | out_product_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      out_product_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      out_product_rsci_bcwt <= 1'b0;
    end
    else begin
      out_product_rsci_bcwt <= ~((~(out_product_rsci_bcwt | out_product_rsci_biwt))
          | out_product_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product_run_out_product_rsci_out_product_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_outer_product_run_out_product_rsci_out_product_wait_ctrl (
  run_wen, out_product_rsci_oswt, out_product_rsci_biwt, out_product_rsci_bdwt, out_product_rsci_bcwt,
      out_product_rsci_irdy, out_product_rsci_ivld_run_sct
);
  input run_wen;
  input out_product_rsci_oswt;
  output out_product_rsci_biwt;
  output out_product_rsci_bdwt;
  input out_product_rsci_bcwt;
  input out_product_rsci_irdy;
  output out_product_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire out_product_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign out_product_rsci_bdwt = out_product_rsci_oswt & run_wen;
  assign out_product_rsci_biwt = out_product_rsci_ogwt & out_product_rsci_irdy;
  assign out_product_rsci_ogwt = out_product_rsci_oswt & (~ out_product_rsci_bcwt);
  assign out_product_rsci_ivld_run_sct = out_product_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product_run_filtered_gradient_rsci_filtered_gradient_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_outer_product_run_filtered_gradient_rsci_filtered_gradient_wait_ctrl
    (
  run_wen, filtered_gradient_rsci_iswt0, filtered_gradient_rsci_irdy_run_sct
);
  input run_wen;
  input filtered_gradient_rsci_iswt0;
  output filtered_gradient_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign filtered_gradient_rsci_irdy_run_sct = filtered_gradient_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product_run_out_product_rsci
// ------------------------------------------------------------------


module OpticalFlow_outer_product_run_out_product_rsci (
  clk, rst, arst_n, out_product_rsc_dat, out_product_rsc_vld, out_product_rsc_rdy,
      run_wen, out_product_rsci_oswt, out_product_rsci_wen_comp, out_product_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [383:0] out_product_rsc_dat;
  output out_product_rsc_vld;
  input out_product_rsc_rdy;
  input run_wen;
  input out_product_rsci_oswt;
  output out_product_rsci_wen_comp;
  input [383:0] out_product_rsci_idat;


  // Interconnect Declarations
  wire out_product_rsci_biwt;
  wire out_product_rsci_bdwt;
  wire out_product_rsci_bcwt;
  wire out_product_rsci_irdy;
  wire out_product_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd384)) out_product_rsci (
      .irdy(out_product_rsci_irdy),
      .ivld(out_product_rsci_ivld_run_sct),
      .idat(out_product_rsci_idat),
      .rdy(out_product_rsc_rdy),
      .vld(out_product_rsc_vld),
      .dat(out_product_rsc_dat)
    );
  OpticalFlow_outer_product_run_out_product_rsci_out_product_wait_ctrl OpticalFlow_outer_product_run_out_product_rsci_out_product_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .out_product_rsci_oswt(out_product_rsci_oswt),
      .out_product_rsci_biwt(out_product_rsci_biwt),
      .out_product_rsci_bdwt(out_product_rsci_bdwt),
      .out_product_rsci_bcwt(out_product_rsci_bcwt),
      .out_product_rsci_irdy(out_product_rsci_irdy),
      .out_product_rsci_ivld_run_sct(out_product_rsci_ivld_run_sct)
    );
  OpticalFlow_outer_product_run_out_product_rsci_out_product_wait_dp OpticalFlow_outer_product_run_out_product_rsci_out_product_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .out_product_rsci_oswt(out_product_rsci_oswt),
      .out_product_rsci_wen_comp(out_product_rsci_wen_comp),
      .out_product_rsci_biwt(out_product_rsci_biwt),
      .out_product_rsci_bdwt(out_product_rsci_bdwt),
      .out_product_rsci_bcwt(out_product_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product_run_filtered_gradient_rsci
// ------------------------------------------------------------------


module OpticalFlow_outer_product_run_filtered_gradient_rsci (
  filtered_gradient_rsc_dat, filtered_gradient_rsc_vld, filtered_gradient_rsc_rdy,
      run_wen, filtered_gradient_rsci_oswt, filtered_gradient_rsci_wen_comp, filtered_gradient_rsci_idat_mxwt
);
  input [95:0] filtered_gradient_rsc_dat;
  input filtered_gradient_rsc_vld;
  output filtered_gradient_rsc_rdy;
  input run_wen;
  input filtered_gradient_rsci_oswt;
  output filtered_gradient_rsci_wen_comp;
  output [95:0] filtered_gradient_rsci_idat_mxwt;


  // Interconnect Declarations
  wire filtered_gradient_rsci_irdy_run_sct;
  wire filtered_gradient_rsci_ivld;
  wire [95:0] filtered_gradient_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd1),
  .width(32'sd96)) filtered_gradient_rsci (
      .rdy(filtered_gradient_rsc_rdy),
      .vld(filtered_gradient_rsc_vld),
      .dat(filtered_gradient_rsc_dat),
      .irdy(filtered_gradient_rsci_irdy_run_sct),
      .ivld(filtered_gradient_rsci_ivld),
      .idat(filtered_gradient_rsci_idat)
    );
  OpticalFlow_outer_product_run_filtered_gradient_rsci_filtered_gradient_wait_ctrl
      OpticalFlow_outer_product_run_filtered_gradient_rsci_filtered_gradient_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .filtered_gradient_rsci_iswt0(filtered_gradient_rsci_oswt),
      .filtered_gradient_rsci_irdy_run_sct(filtered_gradient_rsci_irdy_run_sct)
    );
  assign filtered_gradient_rsci_idat_mxwt = filtered_gradient_rsci_idat;
  assign filtered_gradient_rsci_wen_comp = (~ filtered_gradient_rsci_oswt) | filtered_gradient_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product_run
// ------------------------------------------------------------------


module OpticalFlow_outer_product_run (
  clk, rst, arst_n, filtered_gradient_rsc_dat, filtered_gradient_rsc_vld, filtered_gradient_rsc_rdy,
      out_product_rsc_dat, out_product_rsc_vld, out_product_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [95:0] filtered_gradient_rsc_dat;
  input filtered_gradient_rsc_vld;
  output filtered_gradient_rsc_rdy;
  output [383:0] out_product_rsc_dat;
  output out_product_rsc_vld;
  input out_product_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire filtered_gradient_rsci_wen_comp;
  wire [95:0] filtered_gradient_rsci_idat_mxwt;
  wire out_product_rsci_wen_comp;
  reg [58:0] out_product_rsci_idat_378_320;
  wire [59:0] nl_out_product_rsci_idat_378_320;
  reg [58:0] out_product_rsci_idat_314_256;
  wire [59:0] nl_out_product_rsci_idat_314_256;
  reg [58:0] out_product_rsci_idat_250_192;
  wire [59:0] nl_out_product_rsci_idat_250_192;
  reg [58:0] out_product_rsci_idat_186_128;
  wire [59:0] nl_out_product_rsci_idat_186_128;
  reg [58:0] out_product_rsci_idat_122_64;
  wire [59:0] nl_out_product_rsci_idat_122_64;
  reg [58:0] out_product_rsci_idat_58_0;
  wire [59:0] nl_out_product_rsci_idat_58_0;
  wire [1:0] fsm_output;
  reg main_stage_0_2;
  wire Outer_product_COLUMN_and_cse;
  reg reg_out_product_rsci_iswt0_cse;
  reg reg_filtered_gradient_rsci_iswt0_cse;
  reg [57:0] Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_58_1_itm_1;
  reg Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_0_itm_1;
  reg [57:0] Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_58_1_itm_1;
  reg Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_0_itm_1;
  reg [57:0] Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_58_1_itm_1;
  reg Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_0_itm_1;
  reg [57:0] Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_58_1_itm_1;
  reg Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_0_itm_1;
  reg [57:0] Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_58_1_itm_1;
  reg Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_0_itm_1;
  reg [57:0] Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_58_1_itm_1;
  reg Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_0_itm_1;
  wire [58:0] Outer_product_COLUMN_Outer_product_COLUMN_sqr_itm_63_5_1;
  wire [58:0] Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_itm_63_5_1;
  wire [58:0] Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_itm_63_5_1;
  wire [58:0] Outer_product_COLUMN_Outer_product_COLUMN_mul_itm_63_5_1;
  wire [58:0] Outer_product_COLUMN_Outer_product_COLUMN_mul_1_itm_63_5_1;
  wire [58:0] Outer_product_COLUMN_Outer_product_COLUMN_mul_2_itm_63_5_1;

  wire[63:0] Outer_product_COLUMN_Outer_product_COLUMN_sqr_nl;
  wire signed [63:0] nl_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sgnd;
  wire[63:0] Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_nl;
  wire signed [63:0] nl_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sgnd;
  wire[63:0] Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_nl;
  wire signed [63:0] nl_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sgnd;
  wire[63:0] Outer_product_COLUMN_Outer_product_COLUMN_mul_nl;
  wire signed [63:0] nl_Outer_product_COLUMN_Outer_product_COLUMN_mul_sgnd;
  wire[63:0] Outer_product_COLUMN_Outer_product_COLUMN_mul_1_nl;
  wire signed [63:0] nl_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sgnd;
  wire[63:0] Outer_product_COLUMN_Outer_product_COLUMN_mul_2_nl;
  wire signed [63:0] nl_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sgnd;

  // Interconnect Declarations for Component Instantiations 
  wire [383:0] nl_OpticalFlow_outer_product_run_out_product_rsci_inst_out_product_rsci_idat;
  assign nl_OpticalFlow_outer_product_run_out_product_rsci_inst_out_product_rsci_idat
      = signext_384_379({out_product_rsci_idat_378_320 , ({{5{out_product_rsci_idat_314_256[58]}},
      out_product_rsci_idat_314_256}) , ({{5{out_product_rsci_idat_250_192[58]}},
      out_product_rsci_idat_250_192}) , ({{5{out_product_rsci_idat_186_128[58]}},
      out_product_rsci_idat_186_128}) , ({{5{out_product_rsci_idat_122_64[58]}},
      out_product_rsci_idat_122_64}) , ({{5{out_product_rsci_idat_58_0[58]}}, out_product_rsci_idat_58_0})});
  OpticalFlow_outer_product_run_filtered_gradient_rsci OpticalFlow_outer_product_run_filtered_gradient_rsci_inst
      (
      .filtered_gradient_rsc_dat(filtered_gradient_rsc_dat),
      .filtered_gradient_rsc_vld(filtered_gradient_rsc_vld),
      .filtered_gradient_rsc_rdy(filtered_gradient_rsc_rdy),
      .run_wen(run_wen),
      .filtered_gradient_rsci_oswt(reg_filtered_gradient_rsci_iswt0_cse),
      .filtered_gradient_rsci_wen_comp(filtered_gradient_rsci_wen_comp),
      .filtered_gradient_rsci_idat_mxwt(filtered_gradient_rsci_idat_mxwt)
    );
  OpticalFlow_outer_product_run_out_product_rsci OpticalFlow_outer_product_run_out_product_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .out_product_rsc_dat(out_product_rsc_dat),
      .out_product_rsc_vld(out_product_rsc_vld),
      .out_product_rsc_rdy(out_product_rsc_rdy),
      .run_wen(run_wen),
      .out_product_rsci_oswt(reg_out_product_rsci_iswt0_cse),
      .out_product_rsci_wen_comp(out_product_rsci_wen_comp),
      .out_product_rsci_idat(nl_OpticalFlow_outer_product_run_out_product_rsci_inst_out_product_rsci_idat[383:0])
    );
  OpticalFlow_outer_product_run_staller OpticalFlow_outer_product_run_staller_inst
      (
      .run_wen(run_wen),
      .filtered_gradient_rsci_wen_comp(filtered_gradient_rsci_wen_comp),
      .out_product_rsci_wen_comp(out_product_rsci_wen_comp)
    );
  OpticalFlow_outer_product_run_run_fsm OpticalFlow_outer_product_run_run_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign Outer_product_COLUMN_and_cse = run_wen & main_stage_0_2;
  assign nl_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sgnd = $signed((filtered_gradient_rsci_idat_mxwt[31:0]))
      * $signed((filtered_gradient_rsci_idat_mxwt[31:0]));
  assign Outer_product_COLUMN_Outer_product_COLUMN_sqr_nl = $unsigned(nl_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sgnd);
  assign Outer_product_COLUMN_Outer_product_COLUMN_sqr_itm_63_5_1 = readslicef_64_59_5(Outer_product_COLUMN_Outer_product_COLUMN_sqr_nl);
  assign nl_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sgnd = $signed((filtered_gradient_rsci_idat_mxwt[63:32]))
      * $signed((filtered_gradient_rsci_idat_mxwt[63:32]));
  assign Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_nl = $unsigned(nl_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sgnd);
  assign Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_itm_63_5_1 = readslicef_64_59_5(Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_nl);
  assign nl_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sgnd = $signed((filtered_gradient_rsci_idat_mxwt[95:64]))
      * $signed((filtered_gradient_rsci_idat_mxwt[95:64]));
  assign Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_nl = $unsigned(nl_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sgnd);
  assign Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_itm_63_5_1 = readslicef_64_59_5(Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_nl);
  assign nl_Outer_product_COLUMN_Outer_product_COLUMN_mul_sgnd = $signed((filtered_gradient_rsci_idat_mxwt[31:0]))
      * $signed((filtered_gradient_rsci_idat_mxwt[63:32]));
  assign Outer_product_COLUMN_Outer_product_COLUMN_mul_nl = $unsigned(nl_Outer_product_COLUMN_Outer_product_COLUMN_mul_sgnd);
  assign Outer_product_COLUMN_Outer_product_COLUMN_mul_itm_63_5_1 = readslicef_64_59_5(Outer_product_COLUMN_Outer_product_COLUMN_mul_nl);
  assign nl_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sgnd = $signed((filtered_gradient_rsci_idat_mxwt[31:0]))
      * $signed((filtered_gradient_rsci_idat_mxwt[95:64]));
  assign Outer_product_COLUMN_Outer_product_COLUMN_mul_1_nl = $unsigned(nl_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sgnd);
  assign Outer_product_COLUMN_Outer_product_COLUMN_mul_1_itm_63_5_1 = readslicef_64_59_5(Outer_product_COLUMN_Outer_product_COLUMN_mul_1_nl);
  assign nl_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sgnd = $signed((filtered_gradient_rsci_idat_mxwt[63:32]))
      * $signed((filtered_gradient_rsci_idat_mxwt[95:64]));
  assign Outer_product_COLUMN_Outer_product_COLUMN_mul_2_nl = $unsigned(nl_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sgnd);
  assign Outer_product_COLUMN_Outer_product_COLUMN_mul_2_itm_63_5_1 = readslicef_64_59_5(Outer_product_COLUMN_Outer_product_COLUMN_mul_2_nl);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      out_product_rsci_idat_58_0 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_122_64 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_186_128 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_250_192 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_314_256 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_378_320 <= 59'b00000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      out_product_rsci_idat_58_0 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_122_64 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_186_128 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_250_192 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_314_256 <= 59'b00000000000000000000000000000000000000000000000000000000000;
      out_product_rsci_idat_378_320 <= 59'b00000000000000000000000000000000000000000000000000000000000;
    end
    else if ( Outer_product_COLUMN_and_cse ) begin
      out_product_rsci_idat_58_0 <= nl_out_product_rsci_idat_58_0[58:0];
      out_product_rsci_idat_122_64 <= nl_out_product_rsci_idat_122_64[58:0];
      out_product_rsci_idat_186_128 <= nl_out_product_rsci_idat_186_128[58:0];
      out_product_rsci_idat_250_192 <= nl_out_product_rsci_idat_250_192[58:0];
      out_product_rsci_idat_314_256 <= nl_out_product_rsci_idat_314_256[58:0];
      out_product_rsci_idat_378_320 <= nl_out_product_rsci_idat_378_320[58:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_out_product_rsci_iswt0_cse <= 1'b0;
      reg_filtered_gradient_rsci_iswt0_cse <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_0_itm_1
          <= 1'b0;
      main_stage_0_2 <= 1'b0;
    end
    else if ( rst ) begin
      reg_out_product_rsci_iswt0_cse <= 1'b0;
      reg_filtered_gradient_rsci_iswt0_cse <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_0_itm_1
          <= 1'b0;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_58_1_itm_1
          <= 58'b0000000000000000000000000000000000000000000000000000000000;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_0_itm_1
          <= 1'b0;
      main_stage_0_2 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_out_product_rsci_iswt0_cse <= main_stage_0_2;
      reg_filtered_gradient_rsci_iswt0_cse <= 1'b1;
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_58_1_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_mul_2_itm_63_5_1[58:1];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_0_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_mul_2_itm_63_5_1[0];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_58_1_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_sqr_itm_63_5_1[58:1];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_0_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_sqr_itm_63_5_1[0];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_58_1_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_mul_1_itm_63_5_1[58:1];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_0_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_mul_1_itm_63_5_1[0];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_58_1_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_itm_63_5_1[58:1];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_0_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_itm_63_5_1[0];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_58_1_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_mul_itm_63_5_1[58:1];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_0_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_mul_itm_63_5_1[0];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_58_1_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_itm_63_5_1[58:1];
      Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_0_itm_1
          <= Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_itm_63_5_1[0];
      main_stage_0_2 <= fsm_output[1];
    end
  end
  assign nl_out_product_rsci_idat_58_0  = conv_s2u_58_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_58_1_itm_1)
      + conv_u2u_1_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_sdt_63_5_0_itm_1);
  assign nl_out_product_rsci_idat_122_64  = conv_s2u_58_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_58_1_itm_1)
      + conv_u2u_1_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_1_sdt_63_5_0_itm_1);
  assign nl_out_product_rsci_idat_186_128  = conv_s2u_58_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_58_1_itm_1)
      + conv_u2u_1_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_sqr_2_sdt_63_5_0_itm_1);
  assign nl_out_product_rsci_idat_250_192  = conv_s2u_58_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_58_1_itm_1)
      + conv_u2u_1_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_sdt_63_5_0_itm_1);
  assign nl_out_product_rsci_idat_314_256  = conv_s2u_58_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_58_1_itm_1)
      + conv_u2u_1_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_1_sdt_63_5_0_itm_1);
  assign nl_out_product_rsci_idat_378_320  = conv_s2u_58_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_58_1_itm_1)
      + conv_u2u_1_59(Outer_product_COLUMN_slc_Outer_product_COLUMN_Outer_product_COLUMN_mul_2_sdt_63_5_0_itm_1);

  function automatic [58:0] readslicef_64_59_5;
    input [63:0] vector;
    reg [63:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_64_59_5 = tmp[58:0];
  end
  endfunction


  function automatic [383:0] signext_384_379;
    input [378:0] vector;
  begin
    signext_384_379= {{5{vector[378]}}, vector};
  end
  endfunction


  function automatic [58:0] conv_s2u_58_59 ;
    input [57:0]  vector ;
  begin
    conv_s2u_58_59 = {vector[57], vector};
  end
  endfunction


  function automatic [58:0] conv_u2u_1_59 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_59 = {{58{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product_struct
// ------------------------------------------------------------------


module OpticalFlow_outer_product_struct (
  clk, rst, arst_n, filtered_gradient_rsc_dat_z, filtered_gradient_rsc_dat_y, filtered_gradient_rsc_dat_x,
      filtered_gradient_rsc_vld, filtered_gradient_rsc_rdy, out_product_rsc_dat_val,
      out_product_rsc_vld, out_product_rsc_rdy, widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] filtered_gradient_rsc_dat_z;
  input [31:0] filtered_gradient_rsc_dat_y;
  input [31:0] filtered_gradient_rsc_dat_x;
  input filtered_gradient_rsc_vld;
  output filtered_gradient_rsc_rdy;
  output [383:0] out_product_rsc_dat_val;
  output out_product_rsc_vld;
  input out_product_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;


  // Interconnect Declarations
  wire [383:0] out_product_rsc_dat;


  // Interconnect Declarations for Component Instantiations 
  wire [95:0] nl_OpticalFlow_outer_product_run_inst_filtered_gradient_rsc_dat;
  assign nl_OpticalFlow_outer_product_run_inst_filtered_gradient_rsc_dat = {filtered_gradient_rsc_dat_z
      , filtered_gradient_rsc_dat_y , filtered_gradient_rsc_dat_x};
  OpticalFlow_outer_product_run OpticalFlow_outer_product_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .filtered_gradient_rsc_dat(nl_OpticalFlow_outer_product_run_inst_filtered_gradient_rsc_dat[95:0]),
      .filtered_gradient_rsc_vld(filtered_gradient_rsc_vld),
      .filtered_gradient_rsc_rdy(filtered_gradient_rsc_rdy),
      .out_product_rsc_dat(out_product_rsc_dat),
      .out_product_rsc_vld(out_product_rsc_vld),
      .out_product_rsc_rdy(out_product_rsc_rdy)
    );
  assign out_product_rsc_dat_val = out_product_rsc_dat;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_outer_product
// ------------------------------------------------------------------


module OpticalFlow_outer_product (
  clk, rst, arst_n, filtered_gradient_rsc_dat, filtered_gradient_rsc_vld, filtered_gradient_rsc_rdy,
      out_product_rsc_dat, out_product_rsc_vld, out_product_rsc_rdy, widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [95:0] filtered_gradient_rsc_dat;
  input filtered_gradient_rsc_vld;
  output filtered_gradient_rsc_rdy;
  output [383:0] out_product_rsc_dat;
  output out_product_rsc_vld;
  input out_product_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;


  // Interconnect Declarations
  wire [383:0] out_product_rsc_dat_val;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_OpticalFlow_outer_product_struct_inst_filtered_gradient_rsc_dat_z;
  assign nl_OpticalFlow_outer_product_struct_inst_filtered_gradient_rsc_dat_z = filtered_gradient_rsc_dat[95:64];
  wire [31:0] nl_OpticalFlow_outer_product_struct_inst_filtered_gradient_rsc_dat_y;
  assign nl_OpticalFlow_outer_product_struct_inst_filtered_gradient_rsc_dat_y = filtered_gradient_rsc_dat[63:32];
  wire [31:0] nl_OpticalFlow_outer_product_struct_inst_filtered_gradient_rsc_dat_x;
  assign nl_OpticalFlow_outer_product_struct_inst_filtered_gradient_rsc_dat_x = filtered_gradient_rsc_dat[31:0];
  OpticalFlow_outer_product_struct OpticalFlow_outer_product_struct_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .filtered_gradient_rsc_dat_z(nl_OpticalFlow_outer_product_struct_inst_filtered_gradient_rsc_dat_z[31:0]),
      .filtered_gradient_rsc_dat_y(nl_OpticalFlow_outer_product_struct_inst_filtered_gradient_rsc_dat_y[31:0]),
      .filtered_gradient_rsc_dat_x(nl_OpticalFlow_outer_product_struct_inst_filtered_gradient_rsc_dat_x[31:0]),
      .filtered_gradient_rsc_vld(filtered_gradient_rsc_vld),
      .filtered_gradient_rsc_rdy(filtered_gradient_rsc_rdy),
      .out_product_rsc_dat_val(out_product_rsc_dat_val),
      .out_product_rsc_vld(out_product_rsc_vld),
      .out_product_rsc_rdy(out_product_rsc_rdy),
      .widthIn(11'b00000000000),
      .heightIn(9'b000000000)
    );
  assign out_product_rsc_dat = out_product_rsc_dat_val;
endmodule




//------> ../OpticalFlow_gradient_weight_x.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Sun Jun 16 21:06:12 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_x_run_staller
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_x_run_staller (
  run_wen, y_filtered_rsci_wen_comp, filtered_gradient_rsci_wen_comp
);
  output run_wen;
  input y_filtered_rsci_wen_comp;
  input filtered_gradient_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = y_filtered_rsci_wen_comp & filtered_gradient_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_filtered_gradient_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_filtered_gradient_wait_dp
    (
  clk, rst, arst_n, filtered_gradient_rsci_oswt, filtered_gradient_rsci_wen_comp,
      filtered_gradient_rsci_biwt, filtered_gradient_rsci_bdwt, filtered_gradient_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input filtered_gradient_rsci_oswt;
  output filtered_gradient_rsci_wen_comp;
  input filtered_gradient_rsci_biwt;
  input filtered_gradient_rsci_bdwt;
  output filtered_gradient_rsci_bcwt;
  reg filtered_gradient_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign filtered_gradient_rsci_wen_comp = (~ filtered_gradient_rsci_oswt) | filtered_gradient_rsci_biwt
      | filtered_gradient_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      filtered_gradient_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      filtered_gradient_rsci_bcwt <= 1'b0;
    end
    else begin
      filtered_gradient_rsci_bcwt <= ~((~(filtered_gradient_rsci_bcwt | filtered_gradient_rsci_biwt))
          | filtered_gradient_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_filtered_gradient_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_filtered_gradient_wait_ctrl
    (
  run_wen, filtered_gradient_rsci_oswt, filtered_gradient_rsci_biwt, filtered_gradient_rsci_bdwt,
      filtered_gradient_rsci_bcwt, filtered_gradient_rsci_irdy, filtered_gradient_rsci_ivld_run_sct
);
  input run_wen;
  input filtered_gradient_rsci_oswt;
  output filtered_gradient_rsci_biwt;
  output filtered_gradient_rsci_bdwt;
  input filtered_gradient_rsci_bcwt;
  input filtered_gradient_rsci_irdy;
  output filtered_gradient_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire filtered_gradient_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign filtered_gradient_rsci_bdwt = filtered_gradient_rsci_oswt & run_wen;
  assign filtered_gradient_rsci_biwt = filtered_gradient_rsci_ogwt & filtered_gradient_rsci_irdy;
  assign filtered_gradient_rsci_ogwt = filtered_gradient_rsci_oswt & (~ filtered_gradient_rsci_bcwt);
  assign filtered_gradient_rsci_ivld_run_sct = filtered_gradient_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_x_run_y_filtered_rsci_y_filtered_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_x_run_y_filtered_rsci_y_filtered_wait_ctrl (
  run_wen, y_filtered_rsci_iswt0, y_filtered_rsci_irdy_run_sct
);
  input run_wen;
  input y_filtered_rsci_iswt0;
  output y_filtered_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign y_filtered_rsci_irdy_run_sct = y_filtered_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci (
  clk, rst, arst_n, filtered_gradient_rsc_dat, filtered_gradient_rsc_vld, filtered_gradient_rsc_rdy,
      run_wen, filtered_gradient_rsci_oswt, filtered_gradient_rsci_wen_comp, filtered_gradient_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [95:0] filtered_gradient_rsc_dat;
  output filtered_gradient_rsc_vld;
  input filtered_gradient_rsc_rdy;
  input run_wen;
  input filtered_gradient_rsci_oswt;
  output filtered_gradient_rsci_wen_comp;
  input [95:0] filtered_gradient_rsci_idat;


  // Interconnect Declarations
  wire filtered_gradient_rsci_biwt;
  wire filtered_gradient_rsci_bdwt;
  wire filtered_gradient_rsci_bcwt;
  wire filtered_gradient_rsci_irdy;
  wire filtered_gradient_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd96)) filtered_gradient_rsci (
      .irdy(filtered_gradient_rsci_irdy),
      .ivld(filtered_gradient_rsci_ivld_run_sct),
      .idat(filtered_gradient_rsci_idat),
      .rdy(filtered_gradient_rsc_rdy),
      .vld(filtered_gradient_rsc_vld),
      .dat(filtered_gradient_rsc_dat)
    );
  OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_filtered_gradient_wait_ctrl
      OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_filtered_gradient_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .filtered_gradient_rsci_oswt(filtered_gradient_rsci_oswt),
      .filtered_gradient_rsci_biwt(filtered_gradient_rsci_biwt),
      .filtered_gradient_rsci_bdwt(filtered_gradient_rsci_bdwt),
      .filtered_gradient_rsci_bcwt(filtered_gradient_rsci_bcwt),
      .filtered_gradient_rsci_irdy(filtered_gradient_rsci_irdy),
      .filtered_gradient_rsci_ivld_run_sct(filtered_gradient_rsci_ivld_run_sct)
    );
  OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_filtered_gradient_wait_dp
      OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_filtered_gradient_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .filtered_gradient_rsci_oswt(filtered_gradient_rsci_oswt),
      .filtered_gradient_rsci_wen_comp(filtered_gradient_rsci_wen_comp),
      .filtered_gradient_rsci_biwt(filtered_gradient_rsci_biwt),
      .filtered_gradient_rsci_bdwt(filtered_gradient_rsci_bdwt),
      .filtered_gradient_rsci_bcwt(filtered_gradient_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_x_run_y_filtered_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_x_run_y_filtered_rsci (
  y_filtered_rsc_dat, y_filtered_rsc_vld, y_filtered_rsc_rdy, run_wen, y_filtered_rsci_oswt,
      y_filtered_rsci_wen_comp, y_filtered_rsci_idat_mxwt
);
  input [95:0] y_filtered_rsc_dat;
  input y_filtered_rsc_vld;
  output y_filtered_rsc_rdy;
  input run_wen;
  input y_filtered_rsci_oswt;
  output y_filtered_rsci_wen_comp;
  output [95:0] y_filtered_rsci_idat_mxwt;


  // Interconnect Declarations
  wire y_filtered_rsci_irdy_run_sct;
  wire y_filtered_rsci_ivld;
  wire [95:0] y_filtered_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd1),
  .width(32'sd96)) y_filtered_rsci (
      .rdy(y_filtered_rsc_rdy),
      .vld(y_filtered_rsc_vld),
      .dat(y_filtered_rsc_dat),
      .irdy(y_filtered_rsci_irdy_run_sct),
      .ivld(y_filtered_rsci_ivld),
      .idat(y_filtered_rsci_idat)
    );
  OpticalFlow_gradient_weight_x_run_y_filtered_rsci_y_filtered_wait_ctrl OpticalFlow_gradient_weight_x_run_y_filtered_rsci_y_filtered_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .y_filtered_rsci_iswt0(y_filtered_rsci_oswt),
      .y_filtered_rsci_irdy_run_sct(y_filtered_rsci_irdy_run_sct)
    );
  assign y_filtered_rsci_idat_mxwt = y_filtered_rsci_idat;
  assign y_filtered_rsci_wen_comp = (~ y_filtered_rsci_oswt) | y_filtered_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_x_run
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_x_run (
  clk, rst, arst_n, y_filtered_rsc_dat, y_filtered_rsc_vld, y_filtered_rsc_rdy, filtered_gradient_rsc_dat,
      filtered_gradient_rsc_vld, filtered_gradient_rsc_rdy, widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [95:0] y_filtered_rsc_dat;
  input y_filtered_rsc_vld;
  output y_filtered_rsc_rdy;
  output [95:0] filtered_gradient_rsc_dat;
  output filtered_gradient_rsc_vld;
  input filtered_gradient_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;


  // Interconnect Declarations
  wire run_wen;
  wire y_filtered_rsci_wen_comp;
  wire [95:0] y_filtered_rsci_idat_mxwt;
  wire filtered_gradient_rsci_wen_comp;
  reg [31:0] filtered_gradient_rsci_idat_95_64;
  reg [31:0] filtered_gradient_rsci_idat_63_32;
  reg [31:0] filtered_gradient_rsci_idat_31_0;
  wire [9:0] operator_9_false_acc_tmp;
  wire [10:0] nl_operator_9_false_acc_tmp;
  wire Gradient_weight_x_COLUMN_if_2_unequal_tmp;
  wire and_dcpl_14;
  wire or_dcpl_6;
  wire Gradient_weight_x_COLUMN_Gradient_weight_x_COLUMN_if_2_nor_svs_1;
  reg [10:0] operator_11_false_acc_sdt_sva_1;
  wire [11:0] nl_operator_11_false_acc_sdt_sva_1;
  reg operator_11_false_slc_operator_11_false_acc_10_svs_1;
  reg Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_2;
  reg main_stage_0_4;
  reg Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_1;
  reg main_stage_0_3;
  reg main_stage_0_2;
  reg exitL_exit_Gradient_weight_x_ROW_sva;
  reg main_stage_0_5;
  reg Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_3;
  reg operator_11_false_1_slc_32_itm_3;
  reg Gradient_weight_x_COLUMN_if_slc_operator_11_false_acc_11_svs_st_1;
  reg [10:0] Gradient_weight_x_COLUMN_x_lpi_1_dfm_1;
  wire exit_Gradient_weight_x_ROW_sva_2_mx0w0;
  reg exit_Gradient_weight_x_ROW_sva_2;
  reg reg_filtered_gradient_rsci_oswt_cse;
  wire Gradient_weight_x_COLUMN_if_1_and_cse;
  reg reg_y_filtered_rsci_oswt_cse;
  wire [31:0] gradient_buf0_z_mux_cse;
  wire [31:0] gradient_buf0_y_mux_cse;
  wire [31:0] gradient_buf0_x_mux_cse;
  reg [31:0] gradient_buf5_x_lpi_1;
  reg [31:0] gradient_buf5_y_lpi_1;
  reg [31:0] gradient_buf5_z_lpi_1;
  reg [31:0] gradient_buf0_x_lpi_1_dfm_1;
  reg [31:0] gradient_buf0_x_lpi_1_dfm_2;
  reg [31:0] gradient_buf0_y_lpi_1_dfm_1;
  reg [31:0] gradient_buf0_y_lpi_1_dfm_2;
  reg [31:0] gradient_buf0_z_lpi_1_dfm_1;
  reg [31:0] gradient_buf0_z_lpi_1_dfm_2;
  reg [31:0] gradient_buf1_x_lpi_1_dfm_1;
  reg [31:0] gradient_buf1_x_lpi_1_dfm_2;
  reg [31:0] gradient_buf1_y_lpi_1_dfm_1;
  reg [31:0] gradient_buf1_y_lpi_1_dfm_2;
  reg [31:0] gradient_buf1_z_lpi_1_dfm_1;
  reg [31:0] gradient_buf1_z_lpi_1_dfm_2;
  reg [31:0] gradient_buf2_x_lpi_1_dfm_1;
  reg [31:0] gradient_buf2_x_lpi_1_dfm_2;
  reg [31:0] gradient_buf2_y_lpi_1_dfm_1;
  reg [31:0] gradient_buf2_y_lpi_1_dfm_2;
  reg [31:0] gradient_buf2_z_lpi_1_dfm_1;
  reg [31:0] gradient_buf2_z_lpi_1_dfm_2;
  reg [31:0] gradient_buf3_x_lpi_1_dfm_1;
  reg [31:0] gradient_buf3_x_lpi_1_dfm_2;
  reg [31:0] gradient_buf3_y_lpi_1_dfm_1;
  reg [31:0] gradient_buf3_y_lpi_1_dfm_2;
  reg [31:0] gradient_buf3_z_lpi_1_dfm_1;
  reg [31:0] gradient_buf3_z_lpi_1_dfm_2;
  reg [31:0] gradient_buf4_x_lpi_1_dfm_1;
  reg [31:0] gradient_buf4_x_lpi_1_dfm_2;
  reg [31:0] gradient_buf4_y_lpi_1_dfm_1;
  reg [31:0] gradient_buf4_y_lpi_1_dfm_2;
  reg [31:0] gradient_buf4_z_lpi_1_dfm_1;
  reg [31:0] gradient_buf4_z_lpi_1_dfm_2;
  reg [8:0] Gradient_weight_x_ROW_y_lpi_1_dfm_1;
  reg [31:0] gradient0_x_lpi_1_dfm_1;
  reg [31:0] gradient0_y_lpi_1_dfm_1;
  reg [31:0] gradient0_z_lpi_1_dfm_1;
  reg [60:0] Gradient_weight_x_COLUMN_if_1_mul_15_itm_1;
  wire signed [61:0] nl_Gradient_weight_x_COLUMN_if_1_mul_15_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_16_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_16_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_18_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_18_itm_1;
  reg [60:0] Gradient_weight_x_COLUMN_if_1_mul_19_itm_1;
  wire signed [61:0] nl_Gradient_weight_x_COLUMN_if_1_mul_19_itm_1;
  reg [62:0] Gradient_weight_x_COLUMN_if_1_acc_25_itm_1;
  wire [64:0] nl_Gradient_weight_x_COLUMN_if_1_acc_25_itm_1;
  reg [61:0] Gradient_weight_x_COLUMN_if_1_mul_17_itm_1;
  wire signed [62:0] nl_Gradient_weight_x_COLUMN_if_1_mul_17_itm_1;
  reg [61:0] Gradient_weight_x_COLUMN_if_1_mul_17_itm_2;
  reg [31:0] Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_17_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_20_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_20_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_14_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_14_itm_1;
  reg [60:0] Gradient_weight_x_COLUMN_if_1_acc_21_itm_1;
  wire [61:0] nl_Gradient_weight_x_COLUMN_if_1_acc_21_itm_1;
  reg [60:0] Gradient_weight_x_COLUMN_if_1_mul_8_itm_1;
  wire signed [61:0] nl_Gradient_weight_x_COLUMN_if_1_mul_8_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_9_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_9_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_11_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_11_itm_1;
  reg [60:0] Gradient_weight_x_COLUMN_if_1_mul_12_itm_1;
  wire signed [61:0] nl_Gradient_weight_x_COLUMN_if_1_mul_12_itm_1;
  reg [62:0] Gradient_weight_x_COLUMN_if_1_acc_31_itm_1;
  wire [64:0] nl_Gradient_weight_x_COLUMN_if_1_acc_31_itm_1;
  reg [61:0] Gradient_weight_x_COLUMN_if_1_mul_10_itm_1;
  wire signed [62:0] nl_Gradient_weight_x_COLUMN_if_1_mul_10_itm_1;
  reg [61:0] Gradient_weight_x_COLUMN_if_1_mul_10_itm_2;
  reg [31:0] Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_16_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_13_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_13_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_7_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_7_itm_1;
  reg [60:0] Gradient_weight_x_COLUMN_if_1_acc_27_itm_1;
  wire [61:0] nl_Gradient_weight_x_COLUMN_if_1_acc_27_itm_1;
  reg [60:0] Gradient_weight_x_COLUMN_if_1_mul_1_itm_1;
  wire signed [61:0] nl_Gradient_weight_x_COLUMN_if_1_mul_1_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_2_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_2_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_4_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_4_itm_1;
  reg [60:0] Gradient_weight_x_COLUMN_if_1_mul_5_itm_1;
  wire signed [61:0] nl_Gradient_weight_x_COLUMN_if_1_mul_5_itm_1;
  reg [62:0] Gradient_weight_x_COLUMN_if_1_acc_37_itm_1;
  wire [64:0] nl_Gradient_weight_x_COLUMN_if_1_acc_37_itm_1;
  reg [61:0] Gradient_weight_x_COLUMN_if_1_mul_3_itm_1;
  wire signed [62:0] nl_Gradient_weight_x_COLUMN_if_1_mul_3_itm_1;
  reg [61:0] Gradient_weight_x_COLUMN_if_1_mul_3_itm_2;
  reg [31:0] Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_15_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_6_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_6_itm_1;
  reg [59:0] Gradient_weight_x_COLUMN_if_1_mul_itm_1;
  wire signed [60:0] nl_Gradient_weight_x_COLUMN_if_1_mul_itm_1;
  reg [60:0] Gradient_weight_x_COLUMN_if_1_acc_33_itm_1;
  wire [61:0] nl_Gradient_weight_x_COLUMN_if_1_acc_33_itm_1;
  reg operator_11_false_1_slc_32_itm_1;
  reg operator_11_false_1_slc_32_itm_2;
  wire exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  wire [10:0] Gradient_weight_x_COLUMN_x_lpi_1_dfm_3;
  wire [31:0] gradient_buf5_z_lpi_1_mx0;
  wire [31:0] gradient_buf5_y_lpi_1_mx0;
  wire [31:0] gradient_buf5_x_lpi_1_mx0;
  wire operator_11_false_acc_itm_11_1;

  wire[62:0] Gradient_weight_x_COLUMN_if_1_acc_19_nl;
  wire[63:0] nl_Gradient_weight_x_COLUMN_if_1_acc_19_nl;
  wire[61:0] Gradient_weight_x_COLUMN_if_1_acc_24_nl;
  wire[62:0] nl_Gradient_weight_x_COLUMN_if_1_acc_24_nl;
  wire Gradient_weight_x_COLUMN_if_1_not_4_nl;
  wire[62:0] Gradient_weight_x_COLUMN_if_1_acc_nl;
  wire[63:0] nl_Gradient_weight_x_COLUMN_if_1_acc_nl;
  wire[61:0] Gradient_weight_x_COLUMN_if_1_acc_36_nl;
  wire[62:0] nl_Gradient_weight_x_COLUMN_if_1_acc_36_nl;
  wire Gradient_weight_x_COLUMN_if_1_not_5_nl;
  wire[62:0] Gradient_weight_x_COLUMN_if_1_acc_18_nl;
  wire[63:0] nl_Gradient_weight_x_COLUMN_if_1_acc_18_nl;
  wire[61:0] Gradient_weight_x_COLUMN_if_1_acc_30_nl;
  wire[62:0] nl_Gradient_weight_x_COLUMN_if_1_acc_30_nl;
  wire Gradient_weight_x_COLUMN_if_1_not_6_nl;
  wire[29:0] Gradient_weight_x_COLUMN_if_1_acc_38_nl;
  wire[30:0] nl_Gradient_weight_x_COLUMN_if_1_acc_38_nl;
  wire[29:0] Gradient_weight_x_COLUMN_if_1_acc_40_nl;
  wire[30:0] nl_Gradient_weight_x_COLUMN_if_1_acc_40_nl;
  wire[29:0] Gradient_weight_x_COLUMN_if_1_acc_39_nl;
  wire[30:0] nl_Gradient_weight_x_COLUMN_if_1_acc_39_nl;
  wire[11:0] Gradient_weight_x_COLUMN_aelse_acc_nl;
  wire[12:0] nl_Gradient_weight_x_COLUMN_aelse_acc_nl;
  wire[8:0] Gradient_weight_x_COLUMN_if_2_mux_nl;
  wire[8:0] Gradient_weight_x_ROW_acc_nl;
  wire[9:0] nl_Gradient_weight_x_ROW_acc_nl;
  wire Gradient_weight_x_ROW_not_52_nl;
  wire[10:0] operator_11_false_acc_nl;
  wire[11:0] nl_operator_11_false_acc_nl;
  wire Gradient_weight_x_ROW_not_50_nl;
  wire Gradient_weight_x_ROW_not_51_nl;
  wire Gradient_weight_x_ROW_not_46_nl;
  wire[11:0] operator_11_false_1_acc_nl;
  wire[12:0] nl_operator_11_false_1_acc_nl;
  wire Gradient_weight_x_ROW_not_53_nl;
  wire Gradient_weight_x_ROW_not_54_nl;
  wire Gradient_weight_x_ROW_not_55_nl;
  wire Gradient_weight_x_ROW_not_56_nl;
  wire Gradient_weight_x_ROW_not_57_nl;
  wire Gradient_weight_x_ROW_not_58_nl;
  wire Gradient_weight_x_ROW_not_59_nl;
  wire Gradient_weight_x_ROW_not_60_nl;
  wire Gradient_weight_x_ROW_not_61_nl;
  wire Gradient_weight_x_ROW_not_62_nl;
  wire Gradient_weight_x_ROW_not_63_nl;
  wire Gradient_weight_x_ROW_not_64_nl;
  wire Gradient_weight_x_ROW_not_65_nl;
  wire Gradient_weight_x_ROW_not_66_nl;
  wire Gradient_weight_x_ROW_not_48_nl;
  wire Gradient_weight_x_COLUMN_if_2_Gradient_weight_x_COLUMN_if_2_and_nl;
  wire Gradient_weight_x_ROW_mux_2_nl;
  wire[10:0] Gradient_weight_x_COLUMN_if_2_mux_1_nl;
  wire[10:0] Gradient_weight_x_COLUMN_acc_1_nl;
  wire[11:0] nl_Gradient_weight_x_COLUMN_acc_1_nl;
  wire Gradient_weight_x_ROW_Gradient_weight_x_ROW_Gradient_weight_x_ROW_Gradient_weight_x_ROW_not_nl;
  wire[11:0] operator_11_false_acc_nl_1;
  wire[12:0] nl_operator_11_false_acc_nl_1;

  // Interconnect Declarations for Component Instantiations 
  wire [95:0] nl_OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_inst_filtered_gradient_rsci_idat;
  assign nl_OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_inst_filtered_gradient_rsci_idat
      = {filtered_gradient_rsci_idat_95_64 , filtered_gradient_rsci_idat_63_32 ,
      filtered_gradient_rsci_idat_31_0};
  OpticalFlow_gradient_weight_x_run_y_filtered_rsci OpticalFlow_gradient_weight_x_run_y_filtered_rsci_inst
      (
      .y_filtered_rsc_dat(y_filtered_rsc_dat),
      .y_filtered_rsc_vld(y_filtered_rsc_vld),
      .y_filtered_rsc_rdy(y_filtered_rsc_rdy),
      .run_wen(run_wen),
      .y_filtered_rsci_oswt(reg_y_filtered_rsci_oswt_cse),
      .y_filtered_rsci_wen_comp(y_filtered_rsci_wen_comp),
      .y_filtered_rsci_idat_mxwt(y_filtered_rsci_idat_mxwt)
    );
  OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .filtered_gradient_rsc_dat(filtered_gradient_rsc_dat),
      .filtered_gradient_rsc_vld(filtered_gradient_rsc_vld),
      .filtered_gradient_rsc_rdy(filtered_gradient_rsc_rdy),
      .run_wen(run_wen),
      .filtered_gradient_rsci_oswt(reg_filtered_gradient_rsci_oswt_cse),
      .filtered_gradient_rsci_wen_comp(filtered_gradient_rsci_wen_comp),
      .filtered_gradient_rsci_idat(nl_OpticalFlow_gradient_weight_x_run_filtered_gradient_rsci_inst_filtered_gradient_rsci_idat[95:0])
    );
  OpticalFlow_gradient_weight_x_run_staller OpticalFlow_gradient_weight_x_run_staller_inst
      (
      .run_wen(run_wen),
      .y_filtered_rsci_wen_comp(y_filtered_rsci_wen_comp),
      .filtered_gradient_rsci_wen_comp(filtered_gradient_rsci_wen_comp)
    );
  assign Gradient_weight_x_COLUMN_if_1_and_cse = run_wen & ((main_stage_0_5 & Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_3)
      | and_dcpl_14);
  assign gradient_buf0_x_mux_cse = MUX_v_32_2_2((y_filtered_rsci_idat_mxwt[31:0]),
      gradient_buf0_x_lpi_1_dfm_1, Gradient_weight_x_COLUMN_if_slc_operator_11_false_acc_11_svs_st_1);
  assign gradient_buf0_y_mux_cse = MUX_v_32_2_2((y_filtered_rsci_idat_mxwt[63:32]),
      gradient_buf0_y_lpi_1_dfm_1, Gradient_weight_x_COLUMN_if_slc_operator_11_false_acc_11_svs_st_1);
  assign gradient_buf0_z_mux_cse = MUX_v_32_2_2((y_filtered_rsci_idat_mxwt[95:64]),
      gradient_buf0_z_lpi_1_dfm_1, Gradient_weight_x_COLUMN_if_slc_operator_11_false_acc_11_svs_st_1);
  assign Gradient_weight_x_COLUMN_if_2_unequal_tmp = Gradient_weight_x_COLUMN_x_lpi_1_dfm_1
      != ({(operator_11_false_acc_sdt_sva_1[9:0]) , (widthIn[0])});
  assign Gradient_weight_x_COLUMN_Gradient_weight_x_COLUMN_if_2_nor_svs_1 = ~(Gradient_weight_x_COLUMN_if_2_unequal_tmp
      | (operator_11_false_acc_sdt_sva_1[10]));
  assign Gradient_weight_x_ROW_mux_2_nl = MUX_s_1_2_2(exit_Gradient_weight_x_ROW_sva_2_mx0w0,
      exit_Gradient_weight_x_ROW_sva_2, or_dcpl_6);
  assign Gradient_weight_x_COLUMN_if_2_Gradient_weight_x_COLUMN_if_2_and_nl = Gradient_weight_x_ROW_mux_2_nl
      & Gradient_weight_x_COLUMN_Gradient_weight_x_COLUMN_if_2_nor_svs_1;
  assign exitL_exit_Gradient_weight_x_ROW_sva_mx0 = MUX_s_1_2_2(exitL_exit_Gradient_weight_x_ROW_sva,
      Gradient_weight_x_COLUMN_if_2_Gradient_weight_x_COLUMN_if_2_and_nl, main_stage_0_2);
  assign nl_Gradient_weight_x_COLUMN_acc_1_nl = Gradient_weight_x_COLUMN_x_lpi_1_dfm_1
      + 11'b00000000001;
  assign Gradient_weight_x_COLUMN_acc_1_nl = nl_Gradient_weight_x_COLUMN_acc_1_nl[10:0];
  assign Gradient_weight_x_COLUMN_if_2_mux_1_nl = MUX_v_11_2_2(Gradient_weight_x_COLUMN_acc_1_nl,
      ({{10{exit_Gradient_weight_x_ROW_sva_2_mx0w0}}, exit_Gradient_weight_x_ROW_sva_2_mx0w0}),
      Gradient_weight_x_COLUMN_Gradient_weight_x_COLUMN_if_2_nor_svs_1);
  assign Gradient_weight_x_ROW_Gradient_weight_x_ROW_Gradient_weight_x_ROW_Gradient_weight_x_ROW_not_nl
      = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_COLUMN_x_lpi_1_dfm_3 = MUX_v_11_2_2(11'b00000000000, Gradient_weight_x_COLUMN_if_2_mux_1_nl,
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_Gradient_weight_x_ROW_Gradient_weight_x_ROW_not_nl);
  assign exit_Gradient_weight_x_ROW_sva_2_mx0w0 = ~((Gradient_weight_x_ROW_y_lpi_1_dfm_1
      != (operator_9_false_acc_tmp[8:0])) | (operator_9_false_acc_tmp[9]));
  assign nl_operator_9_false_acc_tmp = conv_u2s_9_10(heightIn) + 10'b1111111111;
  assign operator_9_false_acc_tmp = nl_operator_9_false_acc_tmp[9:0];
  assign nl_operator_11_false_acc_nl_1 = ({1'b1 , widthIn}) + conv_u2s_11_12(~ Gradient_weight_x_COLUMN_x_lpi_1_dfm_3);
  assign operator_11_false_acc_nl_1 = nl_operator_11_false_acc_nl_1[11:0];
  assign operator_11_false_acc_itm_11_1 = readslicef_12_1_11(operator_11_false_acc_nl_1);
  assign gradient_buf5_z_lpi_1_mx0 = MUX_v_32_2_2(gradient_buf5_z_lpi_1, gradient_buf4_z_lpi_1_dfm_2,
      main_stage_0_3);
  assign gradient_buf5_y_lpi_1_mx0 = MUX_v_32_2_2(gradient_buf5_y_lpi_1, gradient_buf4_y_lpi_1_dfm_2,
      main_stage_0_3);
  assign gradient_buf5_x_lpi_1_mx0 = MUX_v_32_2_2(gradient_buf5_x_lpi_1, gradient_buf4_x_lpi_1_dfm_2,
      main_stage_0_3);
  assign and_dcpl_14 = main_stage_0_5 & (~ operator_11_false_1_slc_32_itm_3) & (~
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_3);
  assign or_dcpl_6 = (operator_11_false_acc_sdt_sva_1[10]) | Gradient_weight_x_COLUMN_if_2_unequal_tmp;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_filtered_gradient_rsci_oswt_cse <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_acc_25_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_17_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_21_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_37_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_3_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_33_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_31_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_10_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_27_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      operator_11_false_1_slc_32_itm_3 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_3 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_2 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_1 <= 1'b0;
      exitL_exit_Gradient_weight_x_ROW_sva <= 1'b1;
      Gradient_weight_x_COLUMN_x_lpi_1_dfm_1 <= 11'b00000000000;
      Gradient_weight_x_ROW_y_lpi_1_dfm_1 <= 9'b000000000;
      operator_11_false_acc_sdt_sva_1 <= 11'b00000000000;
      operator_11_false_slc_operator_11_false_acc_10_svs_1 <= 1'b0;
      Gradient_weight_x_COLUMN_if_slc_operator_11_false_acc_11_svs_st_1 <= 1'b0;
      reg_y_filtered_rsci_oswt_cse <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_mul_6_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_1_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_2_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_4_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_5_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_13_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_7_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_8_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_9_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_11_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_12_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_20_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_14_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_15_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_16_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_18_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_19_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      operator_11_false_1_slc_32_itm_2 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_mul_3_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_10_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_17_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      gradient0_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_15_itm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf4_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf3_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf1_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf0_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient0_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_16_itm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf4_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf3_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf1_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf0_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient0_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_17_itm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf4_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf3_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf1_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf0_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      operator_11_false_1_slc_32_itm_1 <= 1'b0;
      gradient_buf5_z_lpi_1 <= 32'b00000000000000000000000000000000;
      gradient_buf5_y_lpi_1 <= 32'b00000000000000000000000000000000;
      gradient_buf5_x_lpi_1 <= 32'b00000000000000000000000000000000;
      gradient_buf4_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf4_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf4_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf3_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf3_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf3_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf1_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf1_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf1_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf0_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf0_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf0_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      reg_filtered_gradient_rsci_oswt_cse <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_acc_25_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_17_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_21_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_37_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_3_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_33_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_31_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_10_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_acc_27_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      operator_11_false_1_slc_32_itm_3 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_3 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_2 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_1 <= 1'b0;
      exitL_exit_Gradient_weight_x_ROW_sva <= 1'b1;
      Gradient_weight_x_COLUMN_x_lpi_1_dfm_1 <= 11'b00000000000;
      Gradient_weight_x_ROW_y_lpi_1_dfm_1 <= 9'b000000000;
      operator_11_false_acc_sdt_sva_1 <= 11'b00000000000;
      operator_11_false_slc_operator_11_false_acc_10_svs_1 <= 1'b0;
      Gradient_weight_x_COLUMN_if_slc_operator_11_false_acc_11_svs_st_1 <= 1'b0;
      reg_y_filtered_rsci_oswt_cse <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_mul_6_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_1_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_2_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_4_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_5_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_13_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_7_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_8_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_9_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_11_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_12_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_20_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_14_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_15_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_16_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_18_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_19_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      operator_11_false_1_slc_32_itm_2 <= 1'b0;
      Gradient_weight_x_COLUMN_if_1_mul_3_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_10_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_x_COLUMN_if_1_mul_17_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      gradient0_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_15_itm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf4_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf3_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf1_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf0_x_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient0_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_16_itm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf4_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf3_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf1_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf0_y_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient0_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_17_itm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf4_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf3_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf1_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      gradient_buf0_z_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      operator_11_false_1_slc_32_itm_1 <= 1'b0;
      gradient_buf5_z_lpi_1 <= 32'b00000000000000000000000000000000;
      gradient_buf5_y_lpi_1 <= 32'b00000000000000000000000000000000;
      gradient_buf5_x_lpi_1 <= 32'b00000000000000000000000000000000;
      gradient_buf4_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf4_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf4_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf3_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf3_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf3_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf2_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf1_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf1_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf1_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf0_z_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf0_y_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      gradient_buf0_x_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_filtered_gradient_rsci_oswt_cse <= (~(operator_11_false_1_slc_32_itm_3
          & (~ Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_3)))
          & main_stage_0_5;
      Gradient_weight_x_COLUMN_if_1_acc_25_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_acc_25_itm_1[62:0];
      Gradient_weight_x_COLUMN_if_1_mul_17_itm_2 <= Gradient_weight_x_COLUMN_if_1_mul_17_itm_1;
      Gradient_weight_x_COLUMN_if_1_acc_21_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_acc_21_itm_1[60:0];
      Gradient_weight_x_COLUMN_if_1_acc_37_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_acc_37_itm_1[62:0];
      Gradient_weight_x_COLUMN_if_1_mul_3_itm_2 <= Gradient_weight_x_COLUMN_if_1_mul_3_itm_1;
      Gradient_weight_x_COLUMN_if_1_acc_33_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_acc_33_itm_1[60:0];
      Gradient_weight_x_COLUMN_if_1_acc_31_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_acc_31_itm_1[62:0];
      Gradient_weight_x_COLUMN_if_1_mul_10_itm_2 <= Gradient_weight_x_COLUMN_if_1_mul_10_itm_1;
      Gradient_weight_x_COLUMN_if_1_acc_27_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_acc_27_itm_1[60:0];
      operator_11_false_1_slc_32_itm_3 <= operator_11_false_1_slc_32_itm_2;
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_3 <= Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_2;
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_2 <= Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_1;
      Gradient_weight_x_COLUMN_if_1_Gradient_weight_x_COLUMN_if_1_and_itm_1 <= (readslicef_12_1_11(Gradient_weight_x_COLUMN_aelse_acc_nl))
          & (~ operator_11_false_slc_operator_11_false_acc_10_svs_1);
      exitL_exit_Gradient_weight_x_ROW_sva <= exitL_exit_Gradient_weight_x_ROW_sva_mx0;
      Gradient_weight_x_COLUMN_x_lpi_1_dfm_1 <= Gradient_weight_x_COLUMN_x_lpi_1_dfm_3;
      Gradient_weight_x_ROW_y_lpi_1_dfm_1 <= MUX_v_9_2_2(9'b000000000, Gradient_weight_x_COLUMN_if_2_mux_nl,
          Gradient_weight_x_ROW_not_52_nl);
      operator_11_false_acc_sdt_sva_1 <= nl_operator_11_false_acc_sdt_sva_1[10:0];
      operator_11_false_slc_operator_11_false_acc_10_svs_1 <= readslicef_11_1_10(operator_11_false_acc_nl);
      Gradient_weight_x_COLUMN_if_slc_operator_11_false_acc_11_svs_st_1 <= operator_11_false_acc_itm_11_1;
      reg_y_filtered_rsci_oswt_cse <= ~ operator_11_false_acc_itm_11_1;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      Gradient_weight_x_COLUMN_if_1_mul_6_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_6_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_1_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_1_itm_1[60:0];
      Gradient_weight_x_COLUMN_if_1_mul_2_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_2_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_4_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_4_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_5_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_5_itm_1[60:0];
      Gradient_weight_x_COLUMN_if_1_mul_13_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_13_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_7_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_7_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_8_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_8_itm_1[60:0];
      Gradient_weight_x_COLUMN_if_1_mul_9_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_9_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_11_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_11_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_12_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_12_itm_1[60:0];
      Gradient_weight_x_COLUMN_if_1_mul_20_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_20_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_14_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_14_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_15_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_15_itm_1[60:0];
      Gradient_weight_x_COLUMN_if_1_mul_16_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_16_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_18_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_18_itm_1[59:0];
      Gradient_weight_x_COLUMN_if_1_mul_19_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_19_itm_1[60:0];
      operator_11_false_1_slc_32_itm_2 <= operator_11_false_1_slc_32_itm_1;
      Gradient_weight_x_COLUMN_if_1_mul_3_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_3_itm_1[61:0];
      Gradient_weight_x_COLUMN_if_1_mul_10_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_10_itm_1[61:0];
      Gradient_weight_x_COLUMN_if_1_mul_17_itm_1 <= nl_Gradient_weight_x_COLUMN_if_1_mul_17_itm_1[61:0];
      gradient0_x_lpi_1_dfm_1 <= gradient_buf0_x_mux_cse;
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_15_itm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf5_x_lpi_1_mx0, Gradient_weight_x_ROW_not_50_nl);
      gradient_buf2_x_lpi_1_dfm_2 <= gradient_buf2_x_lpi_1_dfm_1;
      gradient_buf4_x_lpi_1_dfm_2 <= gradient_buf4_x_lpi_1_dfm_1;
      gradient_buf3_x_lpi_1_dfm_2 <= gradient_buf3_x_lpi_1_dfm_1;
      gradient_buf1_x_lpi_1_dfm_2 <= gradient_buf1_x_lpi_1_dfm_1;
      gradient_buf0_x_lpi_1_dfm_2 <= gradient_buf0_x_lpi_1_dfm_1;
      gradient0_y_lpi_1_dfm_1 <= gradient_buf0_y_mux_cse;
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_16_itm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf5_y_lpi_1_mx0, Gradient_weight_x_ROW_not_51_nl);
      gradient_buf2_y_lpi_1_dfm_2 <= gradient_buf2_y_lpi_1_dfm_1;
      gradient_buf4_y_lpi_1_dfm_2 <= gradient_buf4_y_lpi_1_dfm_1;
      gradient_buf3_y_lpi_1_dfm_2 <= gradient_buf3_y_lpi_1_dfm_1;
      gradient_buf1_y_lpi_1_dfm_2 <= gradient_buf1_y_lpi_1_dfm_1;
      gradient_buf0_y_lpi_1_dfm_2 <= gradient_buf0_y_lpi_1_dfm_1;
      gradient0_z_lpi_1_dfm_1 <= gradient_buf0_z_mux_cse;
      Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_17_itm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf5_z_lpi_1_mx0, Gradient_weight_x_ROW_not_46_nl);
      gradient_buf2_z_lpi_1_dfm_2 <= gradient_buf2_z_lpi_1_dfm_1;
      gradient_buf4_z_lpi_1_dfm_2 <= gradient_buf4_z_lpi_1_dfm_1;
      gradient_buf3_z_lpi_1_dfm_2 <= gradient_buf3_z_lpi_1_dfm_1;
      gradient_buf1_z_lpi_1_dfm_2 <= gradient_buf1_z_lpi_1_dfm_1;
      gradient_buf0_z_lpi_1_dfm_2 <= gradient_buf0_z_lpi_1_dfm_1;
      operator_11_false_1_slc_32_itm_1 <= readslicef_12_1_11(operator_11_false_1_acc_nl);
      gradient_buf5_z_lpi_1 <= gradient_buf5_z_lpi_1_mx0;
      gradient_buf5_y_lpi_1 <= gradient_buf5_y_lpi_1_mx0;
      gradient_buf5_x_lpi_1 <= gradient_buf5_x_lpi_1_mx0;
      gradient_buf4_z_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf3_z_lpi_1_dfm_1, Gradient_weight_x_ROW_not_53_nl);
      gradient_buf4_y_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf3_y_lpi_1_dfm_1, Gradient_weight_x_ROW_not_54_nl);
      gradient_buf4_x_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf3_x_lpi_1_dfm_1, Gradient_weight_x_ROW_not_55_nl);
      gradient_buf3_z_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf2_z_lpi_1_dfm_1, Gradient_weight_x_ROW_not_56_nl);
      gradient_buf3_y_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf2_y_lpi_1_dfm_1, Gradient_weight_x_ROW_not_57_nl);
      gradient_buf3_x_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf2_x_lpi_1_dfm_1, Gradient_weight_x_ROW_not_58_nl);
      gradient_buf2_z_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf1_z_lpi_1_dfm_1, Gradient_weight_x_ROW_not_59_nl);
      gradient_buf2_y_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf1_y_lpi_1_dfm_1, Gradient_weight_x_ROW_not_60_nl);
      gradient_buf2_x_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf1_x_lpi_1_dfm_1, Gradient_weight_x_ROW_not_61_nl);
      gradient_buf1_z_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf0_z_lpi_1_dfm_1, Gradient_weight_x_ROW_not_62_nl);
      gradient_buf1_y_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf0_y_lpi_1_dfm_1, Gradient_weight_x_ROW_not_63_nl);
      gradient_buf1_x_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf0_x_lpi_1_dfm_1, Gradient_weight_x_ROW_not_64_nl);
      gradient_buf0_z_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf0_z_mux_cse, Gradient_weight_x_ROW_not_65_nl);
      gradient_buf0_y_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf0_y_mux_cse, Gradient_weight_x_ROW_not_66_nl);
      gradient_buf0_x_lpi_1_dfm_1 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          gradient_buf0_x_mux_cse, Gradient_weight_x_ROW_not_48_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      filtered_gradient_rsci_idat_95_64 <= 32'b00000000000000000000000000000000;
      filtered_gradient_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
      filtered_gradient_rsci_idat_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      filtered_gradient_rsci_idat_95_64 <= 32'b00000000000000000000000000000000;
      filtered_gradient_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
      filtered_gradient_rsci_idat_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( Gradient_weight_x_COLUMN_if_1_and_cse ) begin
      filtered_gradient_rsci_idat_95_64 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (readslicef_63_32_31(Gradient_weight_x_COLUMN_if_1_acc_19_nl)), Gradient_weight_x_COLUMN_if_1_not_4_nl);
      filtered_gradient_rsci_idat_31_0 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (readslicef_63_32_31(Gradient_weight_x_COLUMN_if_1_acc_nl)), Gradient_weight_x_COLUMN_if_1_not_5_nl);
      filtered_gradient_rsci_idat_63_32 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (readslicef_63_32_31(Gradient_weight_x_COLUMN_if_1_acc_18_nl)), Gradient_weight_x_COLUMN_if_1_not_6_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exit_Gradient_weight_x_ROW_sva_2 <= 1'b0;
    end
    else if ( rst ) begin
      exit_Gradient_weight_x_ROW_sva_2 <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_6 | (~ main_stage_0_2))) ) begin
      exit_Gradient_weight_x_ROW_sva_2 <= exit_Gradient_weight_x_ROW_sva_2_mx0w0;
    end
  end
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_25_itm_1  = conv_s2s_61_63(Gradient_weight_x_COLUMN_if_1_mul_15_itm_1)
      + conv_s2s_61_63({Gradient_weight_x_COLUMN_if_1_mul_16_itm_1 , 1'b0}) + conv_s2s_61_63({Gradient_weight_x_COLUMN_if_1_mul_18_itm_1
      , 1'b0}) + conv_s2s_61_63(Gradient_weight_x_COLUMN_if_1_mul_19_itm_1);
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_38_nl = (Gradient_weight_x_COLUMN_if_1_mul_20_itm_1[59:30])
      + 30'b000000000000000000000000000001;
  assign Gradient_weight_x_COLUMN_if_1_acc_38_nl = nl_Gradient_weight_x_COLUMN_if_1_acc_38_nl[29:0];
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_21_itm_1  = conv_s2s_60_61({Gradient_weight_x_COLUMN_if_1_acc_38_nl
      , (Gradient_weight_x_COLUMN_if_1_mul_20_itm_1[29:0])}) + conv_s2s_60_61(Gradient_weight_x_COLUMN_if_1_mul_14_itm_1);
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_37_itm_1  = conv_s2s_61_63(Gradient_weight_x_COLUMN_if_1_mul_1_itm_1)
      + conv_s2s_61_63({Gradient_weight_x_COLUMN_if_1_mul_2_itm_1 , 1'b0}) + conv_s2s_61_63({Gradient_weight_x_COLUMN_if_1_mul_4_itm_1
      , 1'b0}) + conv_s2s_61_63(Gradient_weight_x_COLUMN_if_1_mul_5_itm_1);
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_40_nl = (Gradient_weight_x_COLUMN_if_1_mul_6_itm_1[59:30])
      + 30'b000000000000000000000000000001;
  assign Gradient_weight_x_COLUMN_if_1_acc_40_nl = nl_Gradient_weight_x_COLUMN_if_1_acc_40_nl[29:0];
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_33_itm_1  = conv_s2s_60_61({Gradient_weight_x_COLUMN_if_1_acc_40_nl
      , (Gradient_weight_x_COLUMN_if_1_mul_6_itm_1[29:0])}) + conv_s2s_60_61(Gradient_weight_x_COLUMN_if_1_mul_itm_1);
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_31_itm_1  = conv_s2s_61_63(Gradient_weight_x_COLUMN_if_1_mul_8_itm_1)
      + conv_s2s_61_63({Gradient_weight_x_COLUMN_if_1_mul_9_itm_1 , 1'b0}) + conv_s2s_61_63({Gradient_weight_x_COLUMN_if_1_mul_11_itm_1
      , 1'b0}) + conv_s2s_61_63(Gradient_weight_x_COLUMN_if_1_mul_12_itm_1);
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_39_nl = (Gradient_weight_x_COLUMN_if_1_mul_13_itm_1[59:30])
      + 30'b000000000000000000000000000001;
  assign Gradient_weight_x_COLUMN_if_1_acc_39_nl = nl_Gradient_weight_x_COLUMN_if_1_acc_39_nl[29:0];
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_27_itm_1  = conv_s2s_60_61({Gradient_weight_x_COLUMN_if_1_acc_39_nl
      , (Gradient_weight_x_COLUMN_if_1_mul_13_itm_1[29:0])}) + conv_s2s_60_61(Gradient_weight_x_COLUMN_if_1_mul_7_itm_1);
  assign nl_Gradient_weight_x_COLUMN_aelse_acc_nl = ({1'b1 , Gradient_weight_x_COLUMN_x_lpi_1_dfm_1})
      + conv_u2u_11_12(~ widthIn) + 12'b000000000001;
  assign Gradient_weight_x_COLUMN_aelse_acc_nl = nl_Gradient_weight_x_COLUMN_aelse_acc_nl[11:0];
  assign nl_Gradient_weight_x_ROW_acc_nl = Gradient_weight_x_ROW_y_lpi_1_dfm_1 +
      9'b000000001;
  assign Gradient_weight_x_ROW_acc_nl = nl_Gradient_weight_x_ROW_acc_nl[8:0];
  assign Gradient_weight_x_COLUMN_if_2_mux_nl = MUX_v_9_2_2(Gradient_weight_x_ROW_acc_nl,
      Gradient_weight_x_ROW_y_lpi_1_dfm_1, or_dcpl_6);
  assign Gradient_weight_x_ROW_not_52_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign nl_operator_11_false_acc_sdt_sva_1  = conv_u2u_10_11(widthIn[10:1]) + 11'b00000000001;
  assign nl_operator_11_false_acc_nl = conv_u2u_10_11(Gradient_weight_x_COLUMN_x_lpi_1_dfm_3[10:1])
      + 11'b11111111101;
  assign operator_11_false_acc_nl = nl_operator_11_false_acc_nl[10:0];
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_6_itm_1  = $signed(Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_15_itm_1)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_itm_1  = $signed(gradient0_x_lpi_1_dfm_1)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_1_itm_1  = $signed(gradient_buf0_x_lpi_1_dfm_2)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_2_itm_1  = $signed(gradient_buf1_x_lpi_1_dfm_2)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_4_itm_1  = $signed(gradient_buf3_x_lpi_1_dfm_2)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_5_itm_1  = $signed(gradient_buf4_x_lpi_1_dfm_2)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_13_itm_1  = $signed(Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_16_itm_1)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_7_itm_1  = $signed(gradient0_y_lpi_1_dfm_1)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_8_itm_1  = $signed(gradient_buf0_y_lpi_1_dfm_2)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_9_itm_1  = $signed(gradient_buf1_y_lpi_1_dfm_2)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_11_itm_1  = $signed(gradient_buf3_y_lpi_1_dfm_2)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_12_itm_1  = $signed(gradient_buf4_y_lpi_1_dfm_2)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_20_itm_1  = $signed(Gradient_weight_x_ROW_Gradient_weight_x_ROW_and_17_itm_1)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_14_itm_1  = $signed(gradient0_z_lpi_1_dfm_1)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_15_itm_1  = $signed(gradient_buf0_z_lpi_1_dfm_2)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_16_itm_1  = $signed(gradient_buf1_z_lpi_1_dfm_2)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_18_itm_1  = $signed(gradient_buf3_z_lpi_1_dfm_2)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_19_itm_1  = $signed(gradient_buf4_z_lpi_1_dfm_2)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_3_itm_1  = $signed(gradient_buf2_x_lpi_1_dfm_2)
      * $signed(31'b0100101001010001000110011100111);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_10_itm_1  = $signed(gradient_buf2_y_lpi_1_dfm_2)
      * $signed(31'b0100101001010001000110011100111);
  assign nl_Gradient_weight_x_COLUMN_if_1_mul_17_itm_1  = $signed(gradient_buf2_z_lpi_1_dfm_2)
      * $signed(31'b0100101001010001000110011100111);
  assign Gradient_weight_x_ROW_not_50_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva;
  assign Gradient_weight_x_ROW_not_51_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva;
  assign Gradient_weight_x_ROW_not_46_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva;
  assign nl_operator_11_false_1_acc_nl = conv_u2s_11_12(Gradient_weight_x_COLUMN_x_lpi_1_dfm_1)
      + 12'b111111111101;
  assign operator_11_false_1_acc_nl = nl_operator_11_false_1_acc_nl[11:0];
  assign Gradient_weight_x_ROW_not_53_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_54_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_55_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_56_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_57_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_58_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_59_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_60_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_61_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_62_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_63_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_64_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_65_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_66_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign Gradient_weight_x_ROW_not_48_nl = ~ exitL_exit_Gradient_weight_x_ROW_sva_mx0;
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_24_nl = Gradient_weight_x_COLUMN_if_1_mul_17_itm_2
      + conv_s2s_61_62(Gradient_weight_x_COLUMN_if_1_acc_21_itm_1);
  assign Gradient_weight_x_COLUMN_if_1_acc_24_nl = nl_Gradient_weight_x_COLUMN_if_1_acc_24_nl[61:0];
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_19_nl = Gradient_weight_x_COLUMN_if_1_acc_25_itm_1
      + conv_s2s_62_63(Gradient_weight_x_COLUMN_if_1_acc_24_nl);
  assign Gradient_weight_x_COLUMN_if_1_acc_19_nl = nl_Gradient_weight_x_COLUMN_if_1_acc_19_nl[62:0];
  assign Gradient_weight_x_COLUMN_if_1_not_4_nl = ~ and_dcpl_14;
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_36_nl = Gradient_weight_x_COLUMN_if_1_mul_3_itm_2
      + conv_s2s_61_62(Gradient_weight_x_COLUMN_if_1_acc_33_itm_1);
  assign Gradient_weight_x_COLUMN_if_1_acc_36_nl = nl_Gradient_weight_x_COLUMN_if_1_acc_36_nl[61:0];
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_nl = Gradient_weight_x_COLUMN_if_1_acc_37_itm_1
      + conv_s2s_62_63(Gradient_weight_x_COLUMN_if_1_acc_36_nl);
  assign Gradient_weight_x_COLUMN_if_1_acc_nl = nl_Gradient_weight_x_COLUMN_if_1_acc_nl[62:0];
  assign Gradient_weight_x_COLUMN_if_1_not_5_nl = ~ and_dcpl_14;
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_30_nl = Gradient_weight_x_COLUMN_if_1_mul_10_itm_2
      + conv_s2s_61_62(Gradient_weight_x_COLUMN_if_1_acc_27_itm_1);
  assign Gradient_weight_x_COLUMN_if_1_acc_30_nl = nl_Gradient_weight_x_COLUMN_if_1_acc_30_nl[61:0];
  assign nl_Gradient_weight_x_COLUMN_if_1_acc_18_nl = Gradient_weight_x_COLUMN_if_1_acc_31_itm_1
      + conv_s2s_62_63(Gradient_weight_x_COLUMN_if_1_acc_30_nl);
  assign Gradient_weight_x_COLUMN_if_1_acc_18_nl = nl_Gradient_weight_x_COLUMN_if_1_acc_18_nl[62:0];
  assign Gradient_weight_x_COLUMN_if_1_not_6_nl = ~ and_dcpl_14;

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction


  function automatic [31:0] readslicef_63_32_31;
    input [62:0] vector;
    reg [62:0] tmp;
  begin
    tmp = vector >> 31;
    readslicef_63_32_31 = tmp[31:0];
  end
  endfunction


  function automatic [60:0] conv_s2s_60_61 ;
    input [59:0]  vector ;
  begin
    conv_s2s_60_61 = {vector[59], vector};
  end
  endfunction


  function automatic [61:0] conv_s2s_61_62 ;
    input [60:0]  vector ;
  begin
    conv_s2s_61_62 = {vector[60], vector};
  end
  endfunction


  function automatic [62:0] conv_s2s_61_63 ;
    input [60:0]  vector ;
  begin
    conv_s2s_61_63 = {{2{vector[60]}}, vector};
  end
  endfunction


  function automatic [62:0] conv_s2s_62_63 ;
    input [61:0]  vector ;
  begin
    conv_s2s_62_63 = {vector[61], vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_x_struct
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_x_struct (
  clk, rst, arst_n, y_filtered_rsc_dat_z, y_filtered_rsc_dat_y, y_filtered_rsc_dat_x,
      y_filtered_rsc_vld, y_filtered_rsc_rdy, filtered_gradient_rsc_dat_z, filtered_gradient_rsc_dat_y,
      filtered_gradient_rsc_dat_x, filtered_gradient_rsc_vld, filtered_gradient_rsc_rdy,
      widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] y_filtered_rsc_dat_z;
  input [31:0] y_filtered_rsc_dat_y;
  input [31:0] y_filtered_rsc_dat_x;
  input y_filtered_rsc_vld;
  output y_filtered_rsc_rdy;
  output [31:0] filtered_gradient_rsc_dat_z;
  output [31:0] filtered_gradient_rsc_dat_y;
  output [31:0] filtered_gradient_rsc_dat_x;
  output filtered_gradient_rsc_vld;
  input filtered_gradient_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;


  // Interconnect Declarations
  wire [95:0] filtered_gradient_rsc_dat;


  // Interconnect Declarations for Component Instantiations 
  wire [95:0] nl_OpticalFlow_gradient_weight_x_run_inst_y_filtered_rsc_dat;
  assign nl_OpticalFlow_gradient_weight_x_run_inst_y_filtered_rsc_dat = {y_filtered_rsc_dat_z
      , y_filtered_rsc_dat_y , y_filtered_rsc_dat_x};
  OpticalFlow_gradient_weight_x_run OpticalFlow_gradient_weight_x_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .y_filtered_rsc_dat(nl_OpticalFlow_gradient_weight_x_run_inst_y_filtered_rsc_dat[95:0]),
      .y_filtered_rsc_vld(y_filtered_rsc_vld),
      .y_filtered_rsc_rdy(y_filtered_rsc_rdy),
      .filtered_gradient_rsc_dat(filtered_gradient_rsc_dat),
      .filtered_gradient_rsc_vld(filtered_gradient_rsc_vld),
      .filtered_gradient_rsc_rdy(filtered_gradient_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn)
    );
  assign filtered_gradient_rsc_dat_x = filtered_gradient_rsc_dat[31:0];
  assign filtered_gradient_rsc_dat_y = filtered_gradient_rsc_dat[63:32];
  assign filtered_gradient_rsc_dat_z = filtered_gradient_rsc_dat[95:64];
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_x
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_x (
  clk, rst, arst_n, y_filtered_rsc_dat, y_filtered_rsc_vld, y_filtered_rsc_rdy, filtered_gradient_rsc_dat,
      filtered_gradient_rsc_vld, filtered_gradient_rsc_rdy, widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [95:0] y_filtered_rsc_dat;
  input y_filtered_rsc_vld;
  output y_filtered_rsc_rdy;
  output [95:0] filtered_gradient_rsc_dat;
  output filtered_gradient_rsc_vld;
  input filtered_gradient_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;


  // Interconnect Declarations
  wire [31:0] filtered_gradient_rsc_dat_z;
  wire [31:0] filtered_gradient_rsc_dat_y;
  wire [31:0] filtered_gradient_rsc_dat_x;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_OpticalFlow_gradient_weight_x_struct_inst_y_filtered_rsc_dat_z;
  assign nl_OpticalFlow_gradient_weight_x_struct_inst_y_filtered_rsc_dat_z = y_filtered_rsc_dat[95:64];
  wire [31:0] nl_OpticalFlow_gradient_weight_x_struct_inst_y_filtered_rsc_dat_y;
  assign nl_OpticalFlow_gradient_weight_x_struct_inst_y_filtered_rsc_dat_y = y_filtered_rsc_dat[63:32];
  wire [31:0] nl_OpticalFlow_gradient_weight_x_struct_inst_y_filtered_rsc_dat_x;
  assign nl_OpticalFlow_gradient_weight_x_struct_inst_y_filtered_rsc_dat_x = y_filtered_rsc_dat[31:0];
  OpticalFlow_gradient_weight_x_struct OpticalFlow_gradient_weight_x_struct_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .y_filtered_rsc_dat_z(nl_OpticalFlow_gradient_weight_x_struct_inst_y_filtered_rsc_dat_z[31:0]),
      .y_filtered_rsc_dat_y(nl_OpticalFlow_gradient_weight_x_struct_inst_y_filtered_rsc_dat_y[31:0]),
      .y_filtered_rsc_dat_x(nl_OpticalFlow_gradient_weight_x_struct_inst_y_filtered_rsc_dat_x[31:0]),
      .y_filtered_rsc_vld(y_filtered_rsc_vld),
      .y_filtered_rsc_rdy(y_filtered_rsc_rdy),
      .filtered_gradient_rsc_dat_z(filtered_gradient_rsc_dat_z),
      .filtered_gradient_rsc_dat_y(filtered_gradient_rsc_dat_y),
      .filtered_gradient_rsc_dat_x(filtered_gradient_rsc_dat_x),
      .filtered_gradient_rsc_vld(filtered_gradient_rsc_vld),
      .filtered_gradient_rsc_rdy(filtered_gradient_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn)
    );
  assign filtered_gradient_rsc_dat = {filtered_gradient_rsc_dat_z , filtered_gradient_rsc_dat_y
      , filtered_gradient_rsc_dat_x};
endmodule




//------> ../OpticalFlow_gradient_weight_y.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Sun Jun 16 21:04:58 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_24_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_24_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_23_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_23_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_22_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_22_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_21_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_21_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_20_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_20_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_19_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_19_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_18_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_18_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_17_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_17_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_16_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_16_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_15_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_15_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_14_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_14_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_13_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_13_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_12_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_12_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_11_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_11_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_10_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_10_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_9_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_9_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_8_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_8_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_7_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_7_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_staller
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_staller (
  run_wen, gradient_x_rsci_wen_comp, gradient_y_rsci_wen_comp, gradient_z_rsci_wen_comp,
      y_filtered_rsci_wen_comp
);
  output run_wen;
  input gradient_x_rsci_wen_comp;
  input gradient_y_rsci_wen_comp;
  input gradient_z_rsci_wen_comp;
  input y_filtered_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = gradient_x_rsci_wen_comp & gradient_y_rsci_wen_comp & gradient_z_rsci_wen_comp
      & y_filtered_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_y_filtered_rsci_y_filtered_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_y_filtered_rsci_y_filtered_wait_dp (
  clk, rst, arst_n, y_filtered_rsci_oswt, y_filtered_rsci_wen_comp, y_filtered_rsci_biwt,
      y_filtered_rsci_bdwt, y_filtered_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input y_filtered_rsci_oswt;
  output y_filtered_rsci_wen_comp;
  input y_filtered_rsci_biwt;
  input y_filtered_rsci_bdwt;
  output y_filtered_rsci_bcwt;
  reg y_filtered_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign y_filtered_rsci_wen_comp = (~ y_filtered_rsci_oswt) | y_filtered_rsci_biwt
      | y_filtered_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      y_filtered_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      y_filtered_rsci_bcwt <= 1'b0;
    end
    else begin
      y_filtered_rsci_bcwt <= ~((~(y_filtered_rsci_bcwt | y_filtered_rsci_biwt))
          | y_filtered_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_y_filtered_rsci_y_filtered_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_y_filtered_rsci_y_filtered_wait_ctrl (
  run_wen, y_filtered_rsci_oswt, y_filtered_rsci_biwt, y_filtered_rsci_bdwt, y_filtered_rsci_bcwt,
      y_filtered_rsci_irdy, y_filtered_rsci_ivld_run_sct
);
  input run_wen;
  input y_filtered_rsci_oswt;
  output y_filtered_rsci_biwt;
  output y_filtered_rsci_bdwt;
  input y_filtered_rsci_bcwt;
  input y_filtered_rsci_irdy;
  output y_filtered_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire y_filtered_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign y_filtered_rsci_bdwt = y_filtered_rsci_oswt & run_wen;
  assign y_filtered_rsci_biwt = y_filtered_rsci_ogwt & y_filtered_rsci_irdy;
  assign y_filtered_rsci_ogwt = y_filtered_rsci_oswt & (~ y_filtered_rsci_bcwt);
  assign y_filtered_rsci_ivld_run_sct = y_filtered_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_gradient_z_rsci_gradient_z_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_gradient_z_rsci_gradient_z_wait_ctrl (
  run_wen, gradient_z_rsci_iswt0, gradient_z_rsci_irdy_run_sct
);
  input run_wen;
  input gradient_z_rsci_iswt0;
  output gradient_z_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign gradient_z_rsci_irdy_run_sct = gradient_z_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_gradient_y_rsci_gradient_y_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_gradient_y_rsci_gradient_y_wait_ctrl (
  run_wen, gradient_y_rsci_iswt0, gradient_y_rsci_irdy_run_sct
);
  input run_wen;
  input gradient_y_rsci_iswt0;
  output gradient_y_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign gradient_y_rsci_irdy_run_sct = gradient_y_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_gradient_x_rsci_gradient_x_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_gradient_x_rsci_gradient_x_wait_ctrl (
  run_wen, gradient_x_rsci_iswt0, gradient_x_rsci_irdy_run_sct
);
  input run_wen;
  input gradient_x_rsci_iswt0;
  output gradient_x_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign gradient_x_rsci_irdy_run_sct = gradient_x_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_y_filtered_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_y_filtered_rsci (
  clk, rst, arst_n, y_filtered_rsc_dat, y_filtered_rsc_vld, y_filtered_rsc_rdy, run_wen,
      y_filtered_rsci_oswt, y_filtered_rsci_wen_comp, y_filtered_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [95:0] y_filtered_rsc_dat;
  output y_filtered_rsc_vld;
  input y_filtered_rsc_rdy;
  input run_wen;
  input y_filtered_rsci_oswt;
  output y_filtered_rsci_wen_comp;
  input [95:0] y_filtered_rsci_idat;


  // Interconnect Declarations
  wire y_filtered_rsci_biwt;
  wire y_filtered_rsci_bdwt;
  wire y_filtered_rsci_bcwt;
  wire y_filtered_rsci_irdy;
  wire y_filtered_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd96)) y_filtered_rsci (
      .irdy(y_filtered_rsci_irdy),
      .ivld(y_filtered_rsci_ivld_run_sct),
      .idat(y_filtered_rsci_idat),
      .rdy(y_filtered_rsc_rdy),
      .vld(y_filtered_rsc_vld),
      .dat(y_filtered_rsc_dat)
    );
  OpticalFlow_gradient_weight_y_run_y_filtered_rsci_y_filtered_wait_ctrl OpticalFlow_gradient_weight_y_run_y_filtered_rsci_y_filtered_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .y_filtered_rsci_oswt(y_filtered_rsci_oswt),
      .y_filtered_rsci_biwt(y_filtered_rsci_biwt),
      .y_filtered_rsci_bdwt(y_filtered_rsci_bdwt),
      .y_filtered_rsci_bcwt(y_filtered_rsci_bcwt),
      .y_filtered_rsci_irdy(y_filtered_rsci_irdy),
      .y_filtered_rsci_ivld_run_sct(y_filtered_rsci_ivld_run_sct)
    );
  OpticalFlow_gradient_weight_y_run_y_filtered_rsci_y_filtered_wait_dp OpticalFlow_gradient_weight_y_run_y_filtered_rsci_y_filtered_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .y_filtered_rsci_oswt(y_filtered_rsci_oswt),
      .y_filtered_rsci_wen_comp(y_filtered_rsci_wen_comp),
      .y_filtered_rsci_biwt(y_filtered_rsci_biwt),
      .y_filtered_rsci_bdwt(y_filtered_rsci_bdwt),
      .y_filtered_rsci_bcwt(y_filtered_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_gradient_z_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_gradient_z_rsci (
  gradient_z_rsc_dat, gradient_z_rsc_vld, gradient_z_rsc_rdy, run_wen, gradient_z_rsci_oswt,
      gradient_z_rsci_wen_comp, gradient_z_rsci_idat_mxwt
);
  input [31:0] gradient_z_rsc_dat;
  input gradient_z_rsc_vld;
  output gradient_z_rsc_rdy;
  input run_wen;
  input gradient_z_rsci_oswt;
  output gradient_z_rsci_wen_comp;
  output [31:0] gradient_z_rsci_idat_mxwt;


  // Interconnect Declarations
  wire gradient_z_rsci_irdy_run_sct;
  wire gradient_z_rsci_ivld;
  wire [31:0] gradient_z_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd3),
  .width(32'sd32)) gradient_z_rsci (
      .rdy(gradient_z_rsc_rdy),
      .vld(gradient_z_rsc_vld),
      .dat(gradient_z_rsc_dat),
      .irdy(gradient_z_rsci_irdy_run_sct),
      .ivld(gradient_z_rsci_ivld),
      .idat(gradient_z_rsci_idat)
    );
  OpticalFlow_gradient_weight_y_run_gradient_z_rsci_gradient_z_wait_ctrl OpticalFlow_gradient_weight_y_run_gradient_z_rsci_gradient_z_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .gradient_z_rsci_iswt0(gradient_z_rsci_oswt),
      .gradient_z_rsci_irdy_run_sct(gradient_z_rsci_irdy_run_sct)
    );
  assign gradient_z_rsci_idat_mxwt = gradient_z_rsci_idat;
  assign gradient_z_rsci_wen_comp = (~ gradient_z_rsci_oswt) | gradient_z_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_gradient_y_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_gradient_y_rsci (
  gradient_y_rsc_dat, gradient_y_rsc_vld, gradient_y_rsc_rdy, run_wen, gradient_y_rsci_oswt,
      gradient_y_rsci_wen_comp, gradient_y_rsci_idat_mxwt
);
  input [31:0] gradient_y_rsc_dat;
  input gradient_y_rsc_vld;
  output gradient_y_rsc_rdy;
  input run_wen;
  input gradient_y_rsci_oswt;
  output gradient_y_rsci_wen_comp;
  output [31:0] gradient_y_rsci_idat_mxwt;


  // Interconnect Declarations
  wire gradient_y_rsci_irdy_run_sct;
  wire gradient_y_rsci_ivld;
  wire [31:0] gradient_y_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd2),
  .width(32'sd32)) gradient_y_rsci (
      .rdy(gradient_y_rsc_rdy),
      .vld(gradient_y_rsc_vld),
      .dat(gradient_y_rsc_dat),
      .irdy(gradient_y_rsci_irdy_run_sct),
      .ivld(gradient_y_rsci_ivld),
      .idat(gradient_y_rsci_idat)
    );
  OpticalFlow_gradient_weight_y_run_gradient_y_rsci_gradient_y_wait_ctrl OpticalFlow_gradient_weight_y_run_gradient_y_rsci_gradient_y_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .gradient_y_rsci_iswt0(gradient_y_rsci_oswt),
      .gradient_y_rsci_irdy_run_sct(gradient_y_rsci_irdy_run_sct)
    );
  assign gradient_y_rsci_idat_mxwt = gradient_y_rsci_idat;
  assign gradient_y_rsci_wen_comp = (~ gradient_y_rsci_oswt) | gradient_y_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run_gradient_x_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run_gradient_x_rsci (
  gradient_x_rsc_dat, gradient_x_rsc_vld, gradient_x_rsc_rdy, run_wen, gradient_x_rsci_oswt,
      gradient_x_rsci_wen_comp, gradient_x_rsci_idat_mxwt
);
  input [31:0] gradient_x_rsc_dat;
  input gradient_x_rsc_vld;
  output gradient_x_rsc_rdy;
  input run_wen;
  input gradient_x_rsci_oswt;
  output gradient_x_rsci_wen_comp;
  output [31:0] gradient_x_rsci_idat_mxwt;


  // Interconnect Declarations
  wire gradient_x_rsci_irdy_run_sct;
  wire gradient_x_rsci_ivld;
  wire [31:0] gradient_x_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd1),
  .width(32'sd32)) gradient_x_rsci (
      .rdy(gradient_x_rsc_rdy),
      .vld(gradient_x_rsc_vld),
      .dat(gradient_x_rsc_dat),
      .irdy(gradient_x_rsci_irdy_run_sct),
      .ivld(gradient_x_rsci_ivld),
      .idat(gradient_x_rsci_idat)
    );
  OpticalFlow_gradient_weight_y_run_gradient_x_rsci_gradient_x_wait_ctrl OpticalFlow_gradient_weight_y_run_gradient_x_rsci_gradient_x_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .gradient_x_rsci_iswt0(gradient_x_rsci_oswt),
      .gradient_x_rsci_irdy_run_sct(gradient_x_rsci_irdy_run_sct)
    );
  assign gradient_x_rsci_idat_mxwt = gradient_x_rsci_idat;
  assign gradient_x_rsci_wen_comp = (~ gradient_x_rsci_oswt) | gradient_x_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_run
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_run (
  clk, rst, arst_n, gradient_x_rsc_dat, gradient_x_rsc_vld, gradient_x_rsc_rdy, gradient_y_rsc_dat,
      gradient_y_rsc_vld, gradient_y_rsc_rdy, gradient_z_rsc_dat, gradient_z_rsc_vld,
      gradient_z_rsc_rdy, y_filtered_rsc_dat, y_filtered_rsc_vld, y_filtered_rsc_rdy,
      widthIn, heightIn, line_buf5_Ix_rsci_clken_d, line_buf5_Ix_rsci_d_d, line_buf5_Ix_rsci_q_d,
      line_buf4_Ix_rsci_d_d, line_buf4_Ix_rsci_q_d, line_buf3_Ix_rsci_d_d, line_buf3_Ix_rsci_q_d,
      line_buf2_Ix_rsci_d_d, line_buf2_Ix_rsci_q_d, line_buf1_Ix_rsci_d_d, line_buf1_Ix_rsci_q_d,
      line_buf0_Ix_rsci_d_d, line_buf0_Ix_rsci_q_d, line_buf5_Iy_rsci_d_d, line_buf5_Iy_rsci_q_d,
      line_buf4_Iy_rsci_d_d, line_buf4_Iy_rsci_q_d, line_buf3_Iy_rsci_d_d, line_buf3_Iy_rsci_q_d,
      line_buf2_Iy_rsci_d_d, line_buf2_Iy_rsci_q_d, line_buf1_Iy_rsci_d_d, line_buf1_Iy_rsci_q_d,
      line_buf0_Iy_rsci_d_d, line_buf0_Iy_rsci_q_d, line_buf5_Iz_rsci_d_d, line_buf5_Iz_rsci_q_d,
      line_buf4_Iz_rsci_d_d, line_buf4_Iz_rsci_q_d, line_buf3_Iz_rsci_d_d, line_buf3_Iz_rsci_q_d,
      line_buf2_Iz_rsci_d_d, line_buf2_Iz_rsci_q_d, line_buf1_Iz_rsci_d_d, line_buf1_Iz_rsci_q_d,
      line_buf0_Iz_rsci_d_d, line_buf0_Iz_rsci_q_d, line_buf5_Ix_rsci_adr_d_pff,
      line_buf5_Ix_rsci_we_d_pff, line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] gradient_x_rsc_dat;
  input gradient_x_rsc_vld;
  output gradient_x_rsc_rdy;
  input [31:0] gradient_y_rsc_dat;
  input gradient_y_rsc_vld;
  output gradient_y_rsc_rdy;
  input [31:0] gradient_z_rsc_dat;
  input gradient_z_rsc_vld;
  output gradient_z_rsc_rdy;
  output [95:0] y_filtered_rsc_dat;
  output y_filtered_rsc_vld;
  input y_filtered_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  output line_buf5_Ix_rsci_clken_d;
  output [63:0] line_buf5_Ix_rsci_d_d;
  input [63:0] line_buf5_Ix_rsci_q_d;
  output [63:0] line_buf4_Ix_rsci_d_d;
  input [63:0] line_buf4_Ix_rsci_q_d;
  output [63:0] line_buf3_Ix_rsci_d_d;
  input [63:0] line_buf3_Ix_rsci_q_d;
  output [63:0] line_buf2_Ix_rsci_d_d;
  input [63:0] line_buf2_Ix_rsci_q_d;
  output [63:0] line_buf1_Ix_rsci_d_d;
  input [63:0] line_buf1_Ix_rsci_q_d;
  output [63:0] line_buf0_Ix_rsci_d_d;
  input [63:0] line_buf0_Ix_rsci_q_d;
  output [63:0] line_buf5_Iy_rsci_d_d;
  input [63:0] line_buf5_Iy_rsci_q_d;
  output [63:0] line_buf4_Iy_rsci_d_d;
  input [63:0] line_buf4_Iy_rsci_q_d;
  output [63:0] line_buf3_Iy_rsci_d_d;
  input [63:0] line_buf3_Iy_rsci_q_d;
  output [63:0] line_buf2_Iy_rsci_d_d;
  input [63:0] line_buf2_Iy_rsci_q_d;
  output [63:0] line_buf1_Iy_rsci_d_d;
  input [63:0] line_buf1_Iy_rsci_q_d;
  output [63:0] line_buf0_Iy_rsci_d_d;
  input [63:0] line_buf0_Iy_rsci_q_d;
  output [63:0] line_buf5_Iz_rsci_d_d;
  input [63:0] line_buf5_Iz_rsci_q_d;
  output [63:0] line_buf4_Iz_rsci_d_d;
  input [63:0] line_buf4_Iz_rsci_q_d;
  output [63:0] line_buf3_Iz_rsci_d_d;
  input [63:0] line_buf3_Iz_rsci_q_d;
  output [63:0] line_buf2_Iz_rsci_d_d;
  input [63:0] line_buf2_Iz_rsci_q_d;
  output [63:0] line_buf1_Iz_rsci_d_d;
  input [63:0] line_buf1_Iz_rsci_q_d;
  output [63:0] line_buf0_Iz_rsci_d_d;
  input [63:0] line_buf0_Iz_rsci_q_d;
  output [8:0] line_buf5_Ix_rsci_adr_d_pff;
  output line_buf5_Ix_rsci_we_d_pff;
  output line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire gradient_x_rsci_wen_comp;
  wire [31:0] gradient_x_rsci_idat_mxwt;
  wire gradient_y_rsci_wen_comp;
  wire [31:0] gradient_y_rsci_idat_mxwt;
  wire gradient_z_rsci_wen_comp;
  wire [31:0] gradient_z_rsci_idat_mxwt;
  wire y_filtered_rsci_wen_comp;
  reg [31:0] y_filtered_rsci_idat_95_64;
  reg [31:0] y_filtered_rsci_idat_63_32;
  reg [31:0] y_filtered_rsci_idat_31_0;
  wire [8:0] operator_9_false_acc_tmp;
  wire [9:0] nl_operator_9_false_acc_tmp;
  wire and_dcpl_21;
  wire or_dcpl_7;
  wire and_dcpl_23;
  reg Gradient_weight_y_COLUMN_Gradient_weight_y_COLUMN_if_4_Gradient_weight_y_COLUMN_if_4_nor_svs_1;
  reg operator_9_false_slc_operator_9_false_acc_8_svs_2;
  wire exitL_exit_Gradient_weight_y_ROW_sva_mx0;
  reg Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_2;
  reg main_stage_0_5;
  reg main_stage_0_2;
  reg [9:0] Gradient_weight_y_COLUMN_x_lpi_1_dfm_1_9_0;
  reg operator_9_false_slc_operator_9_false_acc_8_svs_st_1;
  reg Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_1;
  reg main_stage_0_4;
  reg main_stage_0_3;
  reg main_stage_0_6;
  reg Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_3;
  reg operator_9_false_1_slc_operator_9_false_1_acc_9_itm_3;
  reg Gradient_weight_y_COLUMN_if_slc_Gradient_weight_y_COLUMN_acc_9_svs_1;
  reg Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0;
  wire [8:0] Gradient_weight_y_ROW_y_lpi_1_dfm_1;
  reg [8:0] Gradient_weight_y_ROW_y_lpi_1_dfm_2;
  wire exit_Gradient_weight_y_ROW_sva_2_mx0w0;
  reg [10:0] Gradient_weight_y_COLUMN_x_sva_2_1;
  wire [11:0] nl_Gradient_weight_y_COLUMN_x_sva_2_1;
  reg reg_y_filtered_rsci_oswt_cse;
  wire Gradient_weight_y_COLUMN_if_3_and_cse;
  wire wrbuf0_Iz_and_cse;
  reg reg_gradient_z_rsci_oswt_cse;
  wire rdbuf5_Ix_and_cse;
  wire rdbuf5_Iz_and_1_cse;
  reg [31:0] wrbuf0_Iz_31_0_lpi_1_dfm_2;
  reg [31:0] wrbuf0_Iy_31_0_lpi_1_dfm_2;
  reg [31:0] wrbuf0_Ix_31_0_lpi_1_dfm_2;
  reg [31:0] Ix0_lpi_1;
  reg [31:0] Iy0_lpi_1;
  reg [31:0] Iz0_lpi_1;
  reg [63:0] rdbuf0_Ix_lpi_1_dfm_1;
  reg [63:0] rdbuf1_Ix_lpi_1_dfm_1;
  reg [63:0] rdbuf2_Ix_lpi_1_dfm_1;
  reg [63:0] rdbuf3_Ix_lpi_1_dfm_1;
  reg [63:0] rdbuf4_Ix_lpi_1_dfm_1;
  reg [63:0] rdbuf0_Iy_lpi_1_dfm_1;
  reg [63:0] rdbuf1_Iy_lpi_1_dfm_1;
  reg [63:0] rdbuf2_Iy_lpi_1_dfm_1;
  reg [63:0] rdbuf3_Iy_lpi_1_dfm_1;
  reg [63:0] rdbuf4_Iy_lpi_1_dfm_1;
  reg [63:0] rdbuf0_Iz_lpi_1_dfm_1;
  reg [63:0] rdbuf1_Iz_lpi_1_dfm_1;
  reg [63:0] rdbuf2_Iz_lpi_1_dfm_1;
  reg [63:0] rdbuf3_Iz_lpi_1_dfm_1;
  reg [63:0] rdbuf4_Iz_lpi_1_dfm_1;
  reg [8:0] Gradient_weight_y_ROW_y_lpi_1_dfm_1_1;
  reg [31:0] Ix0_lpi_1_dfm_1_1;
  reg [31:0] Ix0_lpi_1_dfm_1_2;
  reg [31:0] Iy0_lpi_1_dfm_1_1;
  reg [31:0] Iy0_lpi_1_dfm_1_2;
  reg [31:0] Iz0_lpi_1_dfm_1_1;
  reg [31:0] Iz0_lpi_1_dfm_1_2;
  reg [31:0] Gradient_weight_y_COLUMN_mux_38_itm_1;
  reg [60:0] Gradient_weight_y_COLUMN_if_3_mul_15_itm_1;
  wire signed [61:0] nl_Gradient_weight_y_COLUMN_if_3_mul_15_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_37_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_16_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_16_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_35_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_18_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_18_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_34_itm_1;
  reg [60:0] Gradient_weight_y_COLUMN_if_3_mul_19_itm_1;
  wire signed [61:0] nl_Gradient_weight_y_COLUMN_if_3_mul_19_itm_1;
  reg [62:0] Gradient_weight_y_COLUMN_if_3_acc_27_itm_1;
  wire [64:0] nl_Gradient_weight_y_COLUMN_if_3_acc_27_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_36_itm_1;
  reg [61:0] Gradient_weight_y_COLUMN_if_3_mul_17_itm_1;
  wire signed [62:0] nl_Gradient_weight_y_COLUMN_if_3_mul_17_itm_1;
  reg [61:0] Gradient_weight_y_COLUMN_if_3_mul_17_itm_2;
  reg [31:0] Gradient_weight_y_COLUMN_mux_33_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_20_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_20_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_14_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_14_itm_1;
  reg [60:0] Gradient_weight_y_COLUMN_if_3_acc_23_itm_1;
  wire [61:0] nl_Gradient_weight_y_COLUMN_if_3_acc_23_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_32_itm_1;
  reg [60:0] Gradient_weight_y_COLUMN_if_3_mul_8_itm_1;
  wire signed [61:0] nl_Gradient_weight_y_COLUMN_if_3_mul_8_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_31_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_9_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_9_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_29_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_11_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_11_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_28_itm_1;
  reg [60:0] Gradient_weight_y_COLUMN_if_3_mul_12_itm_1;
  wire signed [61:0] nl_Gradient_weight_y_COLUMN_if_3_mul_12_itm_1;
  reg [62:0] Gradient_weight_y_COLUMN_if_3_acc_33_itm_1;
  wire [64:0] nl_Gradient_weight_y_COLUMN_if_3_acc_33_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_30_itm_1;
  reg [61:0] Gradient_weight_y_COLUMN_if_3_mul_10_itm_1;
  wire signed [62:0] nl_Gradient_weight_y_COLUMN_if_3_mul_10_itm_1;
  reg [61:0] Gradient_weight_y_COLUMN_if_3_mul_10_itm_2;
  reg [31:0] Gradient_weight_y_COLUMN_mux_27_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_13_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_13_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_7_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_7_itm_1;
  reg [60:0] Gradient_weight_y_COLUMN_if_3_acc_29_itm_1;
  wire [61:0] nl_Gradient_weight_y_COLUMN_if_3_acc_29_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_26_itm_1;
  reg [60:0] Gradient_weight_y_COLUMN_if_3_mul_1_itm_1;
  wire signed [61:0] nl_Gradient_weight_y_COLUMN_if_3_mul_1_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_25_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_2_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_2_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_23_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_4_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_4_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_22_itm_1;
  reg [60:0] Gradient_weight_y_COLUMN_if_3_mul_5_itm_1;
  wire signed [61:0] nl_Gradient_weight_y_COLUMN_if_3_mul_5_itm_1;
  reg [62:0] Gradient_weight_y_COLUMN_if_3_acc_39_itm_1;
  wire [64:0] nl_Gradient_weight_y_COLUMN_if_3_acc_39_itm_1;
  reg [31:0] Gradient_weight_y_COLUMN_mux_24_itm_1;
  reg [61:0] Gradient_weight_y_COLUMN_if_3_mul_3_itm_1;
  wire signed [62:0] nl_Gradient_weight_y_COLUMN_if_3_mul_3_itm_1;
  reg [61:0] Gradient_weight_y_COLUMN_if_3_mul_3_itm_2;
  reg [31:0] Gradient_weight_y_COLUMN_mux_21_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_6_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_6_itm_1;
  reg [59:0] Gradient_weight_y_COLUMN_if_3_mul_itm_1;
  wire signed [60:0] nl_Gradient_weight_y_COLUMN_if_3_mul_itm_1;
  reg [60:0] Gradient_weight_y_COLUMN_if_3_acc_35_itm_1;
  wire [61:0] nl_Gradient_weight_y_COLUMN_if_3_acc_35_itm_1;
  reg operator_9_false_1_slc_operator_9_false_1_acc_9_itm_1;
  reg operator_9_false_1_slc_operator_9_false_1_acc_9_itm_2;
  reg [31:0] rdbuf5_Ix_lpi_1_63_32;
  reg [31:0] rdbuf5_Iy_lpi_1_63_32;
  reg [31:0] rdbuf5_Iz_lpi_1_63_32;
  reg [31:0] rdbuf5_Ix_lpi_1_dfm_1_63_32;
  reg [31:0] rdbuf5_Iy_lpi_1_dfm_1_63_32;
  reg [31:0] rdbuf5_Iz_lpi_1_dfm_1_63_32;
  reg [31:0] rdbuf0_Ix_lpi_1_63_32;
  reg [31:0] rdbuf1_Ix_lpi_1_63_32;
  reg [31:0] rdbuf2_Ix_lpi_1_63_32;
  reg [31:0] rdbuf3_Ix_lpi_1_63_32;
  reg [31:0] rdbuf4_Ix_lpi_1_63_32;
  reg [31:0] rdbuf0_Iy_lpi_1_63_32;
  reg [31:0] rdbuf1_Iy_lpi_1_63_32;
  reg [31:0] rdbuf2_Iy_lpi_1_63_32;
  reg [31:0] rdbuf3_Iy_lpi_1_63_32;
  reg [31:0] rdbuf4_Iy_lpi_1_63_32;
  reg [31:0] rdbuf0_Iz_lpi_1_63_32;
  reg [31:0] rdbuf1_Iz_lpi_1_63_32;
  reg [31:0] rdbuf2_Iz_lpi_1_63_32;
  reg [31:0] rdbuf3_Iz_lpi_1_63_32;
  reg [31:0] rdbuf4_Iz_lpi_1_63_32;
  wire [31:0] Iz0_lpi_1_mx0;
  wire [31:0] Iy0_lpi_1_mx0;
  wire [31:0] Ix0_lpi_1_mx0;
  wire [10:0] Gradient_weight_y_COLUMN_x_lpi_1_dfm_2;
  wire [11:0] operator_11_false_acc_psp_sva_1;
  wire [12:0] nl_operator_11_false_acc_psp_sva_1;
  wire [63:0] rdbuf3_Iz_lpi_1_dfm_3;
  wire [63:0] rdbuf2_Ix_lpi_1_dfm_3;
  wire [63:0] rdbuf0_Iy_lpi_1_dfm_3;
  wire [63:0] rdbuf3_Ix_lpi_1_dfm_3;
  wire [31:0] wrbuf0_Iy_31_0_lpi_1_dfm_4;
  wire [63:0] rdbuf4_Ix_lpi_1_dfm_3;
  wire [63:0] rdbuf2_Iy_lpi_1_dfm_3;
  wire [63:0] rdbuf0_Iz_lpi_1_dfm_3;
  wire [63:0] rdbuf4_Iy_lpi_1_dfm_3;
  wire [31:0] wrbuf0_Ix_31_0_lpi_1_dfm_4;
  wire [63:0] rdbuf0_Ix_lpi_1_dfm_3;
  wire [31:0] wrbuf0_Iz_31_0_lpi_1_dfm_4;
  wire [63:0] rdbuf1_Iy_lpi_1_dfm_3;
  wire [63:0] rdbuf1_Ix_lpi_1_dfm_3;
  wire [63:0] rdbuf2_Iz_lpi_1_dfm_3;
  wire [63:0] rdbuf4_Iz_lpi_1_dfm_3;
  wire [63:0] rdbuf3_Iy_lpi_1_dfm_3;
  wire [63:0] rdbuf1_Iz_lpi_1_dfm_3;
  wire operator_9_false_acc_itm_9_1;

  wire[62:0] Gradient_weight_y_COLUMN_if_3_acc_21_nl;
  wire[63:0] nl_Gradient_weight_y_COLUMN_if_3_acc_21_nl;
  wire[61:0] Gradient_weight_y_COLUMN_if_3_acc_26_nl;
  wire[62:0] nl_Gradient_weight_y_COLUMN_if_3_acc_26_nl;
  wire Gradient_weight_y_COLUMN_if_3_not_3_nl;
  wire[62:0] Gradient_weight_y_COLUMN_if_3_acc_nl;
  wire[63:0] nl_Gradient_weight_y_COLUMN_if_3_acc_nl;
  wire[61:0] Gradient_weight_y_COLUMN_if_3_acc_38_nl;
  wire[62:0] nl_Gradient_weight_y_COLUMN_if_3_acc_38_nl;
  wire Gradient_weight_y_COLUMN_if_3_not_4_nl;
  wire[62:0] Gradient_weight_y_COLUMN_if_3_acc_20_nl;
  wire[63:0] nl_Gradient_weight_y_COLUMN_if_3_acc_20_nl;
  wire[61:0] Gradient_weight_y_COLUMN_if_3_acc_32_nl;
  wire[62:0] nl_Gradient_weight_y_COLUMN_if_3_acc_32_nl;
  wire Gradient_weight_y_COLUMN_if_3_not_5_nl;
  wire[29:0] Gradient_weight_y_COLUMN_if_3_acc_40_nl;
  wire[30:0] nl_Gradient_weight_y_COLUMN_if_3_acc_40_nl;
  wire[29:0] Gradient_weight_y_COLUMN_if_3_acc_42_nl;
  wire[30:0] nl_Gradient_weight_y_COLUMN_if_3_acc_42_nl;
  wire[29:0] Gradient_weight_y_COLUMN_if_3_acc_41_nl;
  wire[30:0] nl_Gradient_weight_y_COLUMN_if_3_acc_41_nl;
  wire[9:0] Gradient_weight_y_COLUMN_aelse_acc_nl;
  wire[10:0] nl_Gradient_weight_y_COLUMN_aelse_acc_nl;
  wire[8:0] operator_9_false_acc_nl;
  wire[9:0] nl_operator_9_false_acc_nl;
  wire[9:0] operator_9_false_1_acc_nl;
  wire[10:0] nl_operator_9_false_1_acc_nl;
  wire[10:0] Gradient_weight_y_COLUMN_if_4_mux_nl;
  wire Gradient_weight_y_ROW_Gradient_weight_y_ROW_Gradient_weight_y_ROW_Gradient_weight_y_ROW_not_nl;
  wire[8:0] Gradient_weight_y_COLUMN_if_4_mux_1_nl;
  wire[8:0] Gradient_weight_y_ROW_acc_nl;
  wire[9:0] nl_Gradient_weight_y_ROW_acc_nl;
  wire Gradient_weight_y_ROW_not_33_nl;
  wire[9:0] operator_9_false_acc_nl_1;
  wire[10:0] nl_operator_9_false_acc_nl_1;

  // Interconnect Declarations for Component Instantiations 
  wire [95:0] nl_OpticalFlow_gradient_weight_y_run_y_filtered_rsci_inst_y_filtered_rsci_idat;
  assign nl_OpticalFlow_gradient_weight_y_run_y_filtered_rsci_inst_y_filtered_rsci_idat
      = {y_filtered_rsci_idat_95_64 , y_filtered_rsci_idat_63_32 , y_filtered_rsci_idat_31_0};
  OpticalFlow_gradient_weight_y_run_gradient_x_rsci OpticalFlow_gradient_weight_y_run_gradient_x_rsci_inst
      (
      .gradient_x_rsc_dat(gradient_x_rsc_dat),
      .gradient_x_rsc_vld(gradient_x_rsc_vld),
      .gradient_x_rsc_rdy(gradient_x_rsc_rdy),
      .run_wen(run_wen),
      .gradient_x_rsci_oswt(reg_gradient_z_rsci_oswt_cse),
      .gradient_x_rsci_wen_comp(gradient_x_rsci_wen_comp),
      .gradient_x_rsci_idat_mxwt(gradient_x_rsci_idat_mxwt)
    );
  OpticalFlow_gradient_weight_y_run_gradient_y_rsci OpticalFlow_gradient_weight_y_run_gradient_y_rsci_inst
      (
      .gradient_y_rsc_dat(gradient_y_rsc_dat),
      .gradient_y_rsc_vld(gradient_y_rsc_vld),
      .gradient_y_rsc_rdy(gradient_y_rsc_rdy),
      .run_wen(run_wen),
      .gradient_y_rsci_oswt(reg_gradient_z_rsci_oswt_cse),
      .gradient_y_rsci_wen_comp(gradient_y_rsci_wen_comp),
      .gradient_y_rsci_idat_mxwt(gradient_y_rsci_idat_mxwt)
    );
  OpticalFlow_gradient_weight_y_run_gradient_z_rsci OpticalFlow_gradient_weight_y_run_gradient_z_rsci_inst
      (
      .gradient_z_rsc_dat(gradient_z_rsc_dat),
      .gradient_z_rsc_vld(gradient_z_rsc_vld),
      .gradient_z_rsc_rdy(gradient_z_rsc_rdy),
      .run_wen(run_wen),
      .gradient_z_rsci_oswt(reg_gradient_z_rsci_oswt_cse),
      .gradient_z_rsci_wen_comp(gradient_z_rsci_wen_comp),
      .gradient_z_rsci_idat_mxwt(gradient_z_rsci_idat_mxwt)
    );
  OpticalFlow_gradient_weight_y_run_y_filtered_rsci OpticalFlow_gradient_weight_y_run_y_filtered_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .y_filtered_rsc_dat(y_filtered_rsc_dat),
      .y_filtered_rsc_vld(y_filtered_rsc_vld),
      .y_filtered_rsc_rdy(y_filtered_rsc_rdy),
      .run_wen(run_wen),
      .y_filtered_rsci_oswt(reg_y_filtered_rsci_oswt_cse),
      .y_filtered_rsci_wen_comp(y_filtered_rsci_wen_comp),
      .y_filtered_rsci_idat(nl_OpticalFlow_gradient_weight_y_run_y_filtered_rsci_inst_y_filtered_rsci_idat[95:0])
    );
  OpticalFlow_gradient_weight_y_run_staller OpticalFlow_gradient_weight_y_run_staller_inst
      (
      .run_wen(run_wen),
      .gradient_x_rsci_wen_comp(gradient_x_rsci_wen_comp),
      .gradient_y_rsci_wen_comp(gradient_y_rsci_wen_comp),
      .gradient_z_rsci_wen_comp(gradient_z_rsci_wen_comp),
      .y_filtered_rsci_wen_comp(y_filtered_rsci_wen_comp)
    );
  assign line_buf5_Ix_rsci_clken_d = run_wen;
  assign Gradient_weight_y_COLUMN_if_3_and_cse = run_wen & ((main_stage_0_6 & Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_3)
      | and_dcpl_21);
  assign rdbuf4_Iz_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf4_Iz_rsci_q_d, rdbuf4_Iz_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf3_Iz_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf3_Iz_rsci_q_d, rdbuf3_Iz_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf2_Iz_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf2_Iz_rsci_q_d, rdbuf2_Iz_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf1_Iz_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf1_Iz_rsci_q_d, rdbuf1_Iz_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf0_Iz_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf0_Iz_rsci_q_d, rdbuf0_Iz_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf4_Iy_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf4_Iy_rsci_q_d, rdbuf4_Iy_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf3_Iy_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf3_Iy_rsci_q_d, rdbuf3_Iy_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf2_Iy_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf2_Iy_rsci_q_d, rdbuf2_Iy_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf1_Iy_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf1_Iy_rsci_q_d, rdbuf1_Iy_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf0_Iy_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf0_Iy_rsci_q_d, rdbuf0_Iy_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf4_Ix_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf4_Ix_rsci_q_d, rdbuf4_Ix_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf3_Ix_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf3_Ix_rsci_q_d, rdbuf3_Ix_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf2_Ix_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf2_Ix_rsci_q_d, rdbuf2_Ix_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf1_Ix_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf1_Ix_rsci_q_d, rdbuf1_Ix_lpi_1_dfm_1,
      or_dcpl_7);
  assign rdbuf0_Ix_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf0_Ix_rsci_q_d, rdbuf0_Ix_lpi_1_dfm_1,
      or_dcpl_7);
  assign wrbuf0_Iz_and_cse = run_wen & (~ (Gradient_weight_y_COLUMN_x_lpi_1_dfm_1_9_0[0]));
  assign wrbuf0_Iz_31_0_lpi_1_dfm_4 = MUX_v_32_2_2(gradient_z_rsci_idat_mxwt, Iz0_lpi_1_mx0,
      Gradient_weight_y_COLUMN_if_slc_Gradient_weight_y_COLUMN_acc_9_svs_1);
  assign wrbuf0_Iy_31_0_lpi_1_dfm_4 = MUX_v_32_2_2(gradient_y_rsci_idat_mxwt, Iy0_lpi_1_mx0,
      Gradient_weight_y_COLUMN_if_slc_Gradient_weight_y_COLUMN_acc_9_svs_1);
  assign wrbuf0_Ix_31_0_lpi_1_dfm_4 = MUX_v_32_2_2(gradient_x_rsci_idat_mxwt, Ix0_lpi_1_mx0,
      Gradient_weight_y_COLUMN_if_slc_Gradient_weight_y_COLUMN_acc_9_svs_1);
  assign rdbuf5_Ix_and_cse = run_wen & main_stage_0_3;
  assign rdbuf5_Iz_and_1_cse = run_wen & (~ or_dcpl_7);
  assign Iz0_lpi_1_mx0 = MUX_v_32_2_2(Iz0_lpi_1, Iz0_lpi_1_dfm_1_1, main_stage_0_3);
  assign Iy0_lpi_1_mx0 = MUX_v_32_2_2(Iy0_lpi_1, Iy0_lpi_1_dfm_1_1, main_stage_0_3);
  assign Ix0_lpi_1_mx0 = MUX_v_32_2_2(Ix0_lpi_1, Ix0_lpi_1_dfm_1_1, main_stage_0_3);
  assign exitL_exit_Gradient_weight_y_ROW_sva_mx0 = ~((~(exit_Gradient_weight_y_ROW_sva_2_mx0w0
      & Gradient_weight_y_COLUMN_Gradient_weight_y_COLUMN_if_4_Gradient_weight_y_COLUMN_if_4_nor_svs_1))
      & main_stage_0_2);
  assign Gradient_weight_y_COLUMN_if_4_mux_nl = MUX_v_11_2_2(Gradient_weight_y_COLUMN_x_sva_2_1,
      ({{10{exit_Gradient_weight_y_ROW_sva_2_mx0w0}}, exit_Gradient_weight_y_ROW_sva_2_mx0w0}),
      Gradient_weight_y_COLUMN_Gradient_weight_y_COLUMN_if_4_Gradient_weight_y_COLUMN_if_4_nor_svs_1);
  assign Gradient_weight_y_ROW_Gradient_weight_y_ROW_Gradient_weight_y_ROW_Gradient_weight_y_ROW_not_nl
      = ~ exitL_exit_Gradient_weight_y_ROW_sva_mx0;
  assign Gradient_weight_y_COLUMN_x_lpi_1_dfm_2 = MUX_v_11_2_2(11'b00000000000, Gradient_weight_y_COLUMN_if_4_mux_nl,
      Gradient_weight_y_ROW_Gradient_weight_y_ROW_Gradient_weight_y_ROW_Gradient_weight_y_ROW_not_nl);
  assign exit_Gradient_weight_y_ROW_sva_2_mx0w0 = ~((Gradient_weight_y_ROW_y_lpi_1_dfm_1_1
      != ({(operator_9_false_acc_tmp[7:0]) , (heightIn[0])})) | (operator_9_false_acc_tmp[8]));
  assign nl_Gradient_weight_y_ROW_acc_nl = Gradient_weight_y_ROW_y_lpi_1_dfm_1_1
      + 9'b000000001;
  assign Gradient_weight_y_ROW_acc_nl = nl_Gradient_weight_y_ROW_acc_nl[8:0];
  assign Gradient_weight_y_COLUMN_if_4_mux_1_nl = MUX_v_9_2_2(Gradient_weight_y_ROW_y_lpi_1_dfm_1_1,
      Gradient_weight_y_ROW_acc_nl, Gradient_weight_y_COLUMN_Gradient_weight_y_COLUMN_if_4_Gradient_weight_y_COLUMN_if_4_nor_svs_1);
  assign Gradient_weight_y_ROW_not_33_nl = ~ exitL_exit_Gradient_weight_y_ROW_sva_mx0;
  assign Gradient_weight_y_ROW_y_lpi_1_dfm_1 = MUX_v_9_2_2(9'b000000000, Gradient_weight_y_COLUMN_if_4_mux_1_nl,
      Gradient_weight_y_ROW_not_33_nl);
  assign nl_operator_9_false_acc_tmp = conv_u2u_8_9(heightIn[8:1]) + 9'b000000001;
  assign operator_9_false_acc_tmp = nl_operator_9_false_acc_tmp[8:0];
  assign nl_operator_9_false_acc_nl_1 = ({1'b1 , heightIn}) + conv_u2s_9_10(~ Gradient_weight_y_ROW_y_lpi_1_dfm_1);
  assign operator_9_false_acc_nl_1 = nl_operator_9_false_acc_nl_1[9:0];
  assign operator_9_false_acc_itm_9_1 = readslicef_10_1_9(operator_9_false_acc_nl_1);
  assign nl_operator_11_false_acc_psp_sva_1 = conv_u2s_11_12(widthIn) + 12'b111111111111;
  assign operator_11_false_acc_psp_sva_1 = nl_operator_11_false_acc_psp_sva_1[11:0];
  assign and_dcpl_21 = main_stage_0_6 & (~ Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_3)
      & (~ operator_9_false_1_slc_operator_9_false_1_acc_9_itm_3);
  assign or_dcpl_7 = (~ main_stage_0_3) | Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0;
  assign and_dcpl_23 = main_stage_0_3 & (~ Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
  assign line_buf5_Ix_rsci_adr_d_pff = Gradient_weight_y_COLUMN_x_lpi_1_dfm_1_9_0[9:1];
  assign line_buf5_Ix_rsci_d_d = rdbuf4_Ix_lpi_1_dfm_3;
  assign line_buf5_Ix_rsci_we_d_pff = (Gradient_weight_y_COLUMN_x_lpi_1_dfm_1_9_0[0])
      & main_stage_0_2;
  assign line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff = ~((Gradient_weight_y_COLUMN_x_lpi_1_dfm_1_9_0[0])
      | (~ main_stage_0_2));
  assign line_buf4_Ix_rsci_d_d = rdbuf3_Ix_lpi_1_dfm_3;
  assign line_buf3_Ix_rsci_d_d = rdbuf2_Ix_lpi_1_dfm_3;
  assign line_buf2_Ix_rsci_d_d = rdbuf1_Ix_lpi_1_dfm_3;
  assign line_buf1_Ix_rsci_d_d = rdbuf0_Ix_lpi_1_dfm_3;
  assign line_buf0_Ix_rsci_d_d = {wrbuf0_Ix_31_0_lpi_1_dfm_4 , wrbuf0_Ix_31_0_lpi_1_dfm_2};
  assign line_buf5_Iy_rsci_d_d = rdbuf4_Iy_lpi_1_dfm_3;
  assign line_buf4_Iy_rsci_d_d = rdbuf3_Iy_lpi_1_dfm_3;
  assign line_buf3_Iy_rsci_d_d = rdbuf2_Iy_lpi_1_dfm_3;
  assign line_buf2_Iy_rsci_d_d = rdbuf1_Iy_lpi_1_dfm_3;
  assign line_buf1_Iy_rsci_d_d = rdbuf0_Iy_lpi_1_dfm_3;
  assign line_buf0_Iy_rsci_d_d = {wrbuf0_Iy_31_0_lpi_1_dfm_4 , wrbuf0_Iy_31_0_lpi_1_dfm_2};
  assign line_buf5_Iz_rsci_d_d = rdbuf4_Iz_lpi_1_dfm_3;
  assign line_buf4_Iz_rsci_d_d = rdbuf3_Iz_lpi_1_dfm_3;
  assign line_buf3_Iz_rsci_d_d = rdbuf2_Iz_lpi_1_dfm_3;
  assign line_buf2_Iz_rsci_d_d = rdbuf1_Iz_lpi_1_dfm_3;
  assign line_buf1_Iz_rsci_d_d = rdbuf0_Iz_lpi_1_dfm_3;
  assign line_buf0_Iz_rsci_d_d = {wrbuf0_Iz_31_0_lpi_1_dfm_4 , wrbuf0_Iz_31_0_lpi_1_dfm_2};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_y_filtered_rsci_oswt_cse <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_acc_27_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_17_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_23_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_39_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_3_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_35_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_33_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_10_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_29_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm_3 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_3 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_2 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_1 <= 1'b0;
      Iz0_lpi_1 <= 32'b00000000000000000000000000000000;
      Iy0_lpi_1 <= 32'b00000000000000000000000000000000;
      Ix0_lpi_1 <= 32'b00000000000000000000000000000000;
      rdbuf4_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf3_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf2_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf1_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf0_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf4_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf3_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf2_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf1_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf0_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf4_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf3_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf2_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf1_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf0_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_ROW_y_lpi_1_dfm_2 <= 9'b000000000;
      Iz0_lpi_1_dfm_1_1 <= 32'b00000000000000000000000000000000;
      Iy0_lpi_1_dfm_1_1 <= 32'b00000000000000000000000000000000;
      Ix0_lpi_1_dfm_1_1 <= 32'b00000000000000000000000000000000;
      operator_9_false_slc_operator_9_false_acc_8_svs_2 <= 1'b0;
      Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0 <= 1'b0;
      Gradient_weight_y_COLUMN_x_lpi_1_dfm_1_9_0 <= 10'b0000000000;
      Gradient_weight_y_COLUMN_Gradient_weight_y_COLUMN_if_4_Gradient_weight_y_COLUMN_if_4_nor_svs_1
          <= 1'b0;
      Gradient_weight_y_ROW_y_lpi_1_dfm_1_1 <= 9'b000000000;
      Gradient_weight_y_COLUMN_x_sva_2_1 <= 11'b00000000000;
      Gradient_weight_y_COLUMN_if_slc_Gradient_weight_y_COLUMN_acc_9_svs_1 <= 1'b0;
      reg_gradient_z_rsci_oswt_cse <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      main_stage_0_6 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_mul_6_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_1_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_2_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_4_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_5_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_13_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_7_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_8_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_9_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_11_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_12_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_20_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_14_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_15_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_16_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_18_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_19_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm_2 <= 1'b0;
      operator_9_false_slc_operator_9_false_acc_8_svs_st_1 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_mul_3_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_10_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_17_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Ix0_lpi_1_dfm_1_2 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_21_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_24_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_22_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_23_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_25_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_26_itm_1 <= 32'b00000000000000000000000000000000;
      Iy0_lpi_1_dfm_1_2 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_27_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_30_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_28_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_29_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_31_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_32_itm_1 <= 32'b00000000000000000000000000000000;
      Iz0_lpi_1_dfm_1_2 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_33_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_36_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_34_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_35_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_37_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_38_itm_1 <= 32'b00000000000000000000000000000000;
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm_1 <= 1'b0;
    end
    else if ( rst ) begin
      reg_y_filtered_rsci_oswt_cse <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_acc_27_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_17_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_23_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_39_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_3_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_35_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_33_itm_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_10_itm_2 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_acc_29_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm_3 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_3 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_2 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_1 <= 1'b0;
      Iz0_lpi_1 <= 32'b00000000000000000000000000000000;
      Iy0_lpi_1 <= 32'b00000000000000000000000000000000;
      Ix0_lpi_1 <= 32'b00000000000000000000000000000000;
      rdbuf4_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf3_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf2_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf1_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf0_Iz_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf4_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf3_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf2_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf1_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf0_Iy_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf4_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf3_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf2_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf1_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf0_Ix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_ROW_y_lpi_1_dfm_2 <= 9'b000000000;
      Iz0_lpi_1_dfm_1_1 <= 32'b00000000000000000000000000000000;
      Iy0_lpi_1_dfm_1_1 <= 32'b00000000000000000000000000000000;
      Ix0_lpi_1_dfm_1_1 <= 32'b00000000000000000000000000000000;
      operator_9_false_slc_operator_9_false_acc_8_svs_2 <= 1'b0;
      Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0 <= 1'b0;
      Gradient_weight_y_COLUMN_x_lpi_1_dfm_1_9_0 <= 10'b0000000000;
      Gradient_weight_y_COLUMN_Gradient_weight_y_COLUMN_if_4_Gradient_weight_y_COLUMN_if_4_nor_svs_1
          <= 1'b0;
      Gradient_weight_y_ROW_y_lpi_1_dfm_1_1 <= 9'b000000000;
      Gradient_weight_y_COLUMN_x_sva_2_1 <= 11'b00000000000;
      Gradient_weight_y_COLUMN_if_slc_Gradient_weight_y_COLUMN_acc_9_svs_1 <= 1'b0;
      reg_gradient_z_rsci_oswt_cse <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      main_stage_0_6 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_mul_6_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_1_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_2_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_4_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_5_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_13_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_7_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_8_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_9_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_11_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_12_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_20_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_14_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_15_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_16_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_18_itm_1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_19_itm_1 <= 61'b0000000000000000000000000000000000000000000000000000000000000;
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm_2 <= 1'b0;
      operator_9_false_slc_operator_9_false_acc_8_svs_st_1 <= 1'b0;
      Gradient_weight_y_COLUMN_if_3_mul_3_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_10_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Gradient_weight_y_COLUMN_if_3_mul_17_itm_1 <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      Ix0_lpi_1_dfm_1_2 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_21_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_24_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_22_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_23_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_25_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_26_itm_1 <= 32'b00000000000000000000000000000000;
      Iy0_lpi_1_dfm_1_2 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_27_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_30_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_28_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_29_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_31_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_32_itm_1 <= 32'b00000000000000000000000000000000;
      Iz0_lpi_1_dfm_1_2 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_33_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_36_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_34_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_35_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_37_itm_1 <= 32'b00000000000000000000000000000000;
      Gradient_weight_y_COLUMN_mux_38_itm_1 <= 32'b00000000000000000000000000000000;
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm_1 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_y_filtered_rsci_oswt_cse <= (~((~ Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_3)
          & operator_9_false_1_slc_operator_9_false_1_acc_9_itm_3)) & main_stage_0_6;
      Gradient_weight_y_COLUMN_if_3_acc_27_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_acc_27_itm_1[62:0];
      Gradient_weight_y_COLUMN_if_3_mul_17_itm_2 <= Gradient_weight_y_COLUMN_if_3_mul_17_itm_1;
      Gradient_weight_y_COLUMN_if_3_acc_23_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_acc_23_itm_1[60:0];
      Gradient_weight_y_COLUMN_if_3_acc_39_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_acc_39_itm_1[62:0];
      Gradient_weight_y_COLUMN_if_3_mul_3_itm_2 <= Gradient_weight_y_COLUMN_if_3_mul_3_itm_1;
      Gradient_weight_y_COLUMN_if_3_acc_35_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_acc_35_itm_1[60:0];
      Gradient_weight_y_COLUMN_if_3_acc_33_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_acc_33_itm_1[62:0];
      Gradient_weight_y_COLUMN_if_3_mul_10_itm_2 <= Gradient_weight_y_COLUMN_if_3_mul_10_itm_1;
      Gradient_weight_y_COLUMN_if_3_acc_29_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_acc_29_itm_1[60:0];
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm_3 <= operator_9_false_1_slc_operator_9_false_1_acc_9_itm_2;
      Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_3 <= Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_2;
      Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_2 <= Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_1;
      Gradient_weight_y_COLUMN_if_3_Gradient_weight_y_COLUMN_if_3_and_itm_1 <= (readslicef_10_1_9(Gradient_weight_y_COLUMN_aelse_acc_nl))
          & (~ operator_9_false_slc_operator_9_false_acc_8_svs_2);
      Iz0_lpi_1 <= Iz0_lpi_1_mx0;
      Iy0_lpi_1 <= Iy0_lpi_1_mx0;
      Ix0_lpi_1 <= Ix0_lpi_1_mx0;
      rdbuf4_Iz_lpi_1_dfm_1 <= rdbuf4_Iz_lpi_1_dfm_3;
      rdbuf3_Iz_lpi_1_dfm_1 <= rdbuf3_Iz_lpi_1_dfm_3;
      rdbuf2_Iz_lpi_1_dfm_1 <= rdbuf2_Iz_lpi_1_dfm_3;
      rdbuf1_Iz_lpi_1_dfm_1 <= rdbuf1_Iz_lpi_1_dfm_3;
      rdbuf0_Iz_lpi_1_dfm_1 <= rdbuf0_Iz_lpi_1_dfm_3;
      rdbuf4_Iy_lpi_1_dfm_1 <= rdbuf4_Iy_lpi_1_dfm_3;
      rdbuf3_Iy_lpi_1_dfm_1 <= rdbuf3_Iy_lpi_1_dfm_3;
      rdbuf2_Iy_lpi_1_dfm_1 <= rdbuf2_Iy_lpi_1_dfm_3;
      rdbuf1_Iy_lpi_1_dfm_1 <= rdbuf1_Iy_lpi_1_dfm_3;
      rdbuf0_Iy_lpi_1_dfm_1 <= rdbuf0_Iy_lpi_1_dfm_3;
      rdbuf4_Ix_lpi_1_dfm_1 <= rdbuf4_Ix_lpi_1_dfm_3;
      rdbuf3_Ix_lpi_1_dfm_1 <= rdbuf3_Ix_lpi_1_dfm_3;
      rdbuf2_Ix_lpi_1_dfm_1 <= rdbuf2_Ix_lpi_1_dfm_3;
      rdbuf1_Ix_lpi_1_dfm_1 <= rdbuf1_Ix_lpi_1_dfm_3;
      rdbuf0_Ix_lpi_1_dfm_1 <= rdbuf0_Ix_lpi_1_dfm_3;
      Gradient_weight_y_ROW_y_lpi_1_dfm_2 <= Gradient_weight_y_ROW_y_lpi_1_dfm_1_1;
      Iz0_lpi_1_dfm_1_1 <= wrbuf0_Iz_31_0_lpi_1_dfm_4;
      Iy0_lpi_1_dfm_1_1 <= wrbuf0_Iy_31_0_lpi_1_dfm_4;
      Ix0_lpi_1_dfm_1_1 <= wrbuf0_Ix_31_0_lpi_1_dfm_4;
      operator_9_false_slc_operator_9_false_acc_8_svs_2 <= operator_9_false_slc_operator_9_false_acc_8_svs_st_1;
      Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0 <= Gradient_weight_y_COLUMN_x_lpi_1_dfm_1_9_0[0];
      Gradient_weight_y_COLUMN_x_lpi_1_dfm_1_9_0 <= Gradient_weight_y_COLUMN_x_lpi_1_dfm_2[9:0];
      Gradient_weight_y_COLUMN_Gradient_weight_y_COLUMN_if_4_Gradient_weight_y_COLUMN_if_4_nor_svs_1
          <= ~((Gradient_weight_y_COLUMN_x_lpi_1_dfm_2 != (operator_11_false_acc_psp_sva_1[10:0]))
          | (operator_11_false_acc_psp_sva_1[11]));
      Gradient_weight_y_ROW_y_lpi_1_dfm_1_1 <= Gradient_weight_y_ROW_y_lpi_1_dfm_1;
      Gradient_weight_y_COLUMN_x_sva_2_1 <= nl_Gradient_weight_y_COLUMN_x_sva_2_1[10:0];
      Gradient_weight_y_COLUMN_if_slc_Gradient_weight_y_COLUMN_acc_9_svs_1 <= operator_9_false_acc_itm_9_1;
      reg_gradient_z_rsci_oswt_cse <= ~ operator_9_false_acc_itm_9_1;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      main_stage_0_6 <= main_stage_0_5;
      Gradient_weight_y_COLUMN_if_3_mul_6_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_6_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_1_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_1_itm_1[60:0];
      Gradient_weight_y_COLUMN_if_3_mul_2_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_2_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_4_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_4_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_5_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_5_itm_1[60:0];
      Gradient_weight_y_COLUMN_if_3_mul_13_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_13_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_7_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_7_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_8_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_8_itm_1[60:0];
      Gradient_weight_y_COLUMN_if_3_mul_9_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_9_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_11_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_11_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_12_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_12_itm_1[60:0];
      Gradient_weight_y_COLUMN_if_3_mul_20_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_20_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_14_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_14_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_15_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_15_itm_1[60:0];
      Gradient_weight_y_COLUMN_if_3_mul_16_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_16_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_18_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_18_itm_1[59:0];
      Gradient_weight_y_COLUMN_if_3_mul_19_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_19_itm_1[60:0];
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm_2 <= operator_9_false_1_slc_operator_9_false_1_acc_9_itm_1;
      operator_9_false_slc_operator_9_false_acc_8_svs_st_1 <= readslicef_9_1_8(operator_9_false_acc_nl);
      Gradient_weight_y_COLUMN_if_3_mul_3_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_3_itm_1[61:0];
      Gradient_weight_y_COLUMN_if_3_mul_10_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_10_itm_1[61:0];
      Gradient_weight_y_COLUMN_if_3_mul_17_itm_1 <= nl_Gradient_weight_y_COLUMN_if_3_mul_17_itm_1[61:0];
      Ix0_lpi_1_dfm_1_2 <= Ix0_lpi_1_dfm_1_1;
      Gradient_weight_y_COLUMN_mux_21_itm_1 <= MUX_v_32_2_2((line_buf5_Ix_rsci_q_d[31:0]),
          rdbuf5_Ix_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_24_itm_1 <= MUX_v_32_2_2((line_buf2_Ix_rsci_q_d[31:0]),
          rdbuf2_Ix_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_22_itm_1 <= MUX_v_32_2_2((line_buf4_Ix_rsci_q_d[31:0]),
          rdbuf4_Ix_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_23_itm_1 <= MUX_v_32_2_2((line_buf3_Ix_rsci_q_d[31:0]),
          rdbuf3_Ix_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_25_itm_1 <= MUX_v_32_2_2((line_buf1_Ix_rsci_q_d[31:0]),
          rdbuf1_Ix_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_26_itm_1 <= MUX_v_32_2_2((line_buf0_Ix_rsci_q_d[31:0]),
          rdbuf0_Ix_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Iy0_lpi_1_dfm_1_2 <= Iy0_lpi_1_dfm_1_1;
      Gradient_weight_y_COLUMN_mux_27_itm_1 <= MUX_v_32_2_2((line_buf5_Iy_rsci_q_d[31:0]),
          rdbuf5_Iy_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_30_itm_1 <= MUX_v_32_2_2((line_buf2_Iy_rsci_q_d[31:0]),
          rdbuf2_Iy_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_28_itm_1 <= MUX_v_32_2_2((line_buf4_Iy_rsci_q_d[31:0]),
          rdbuf4_Iy_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_29_itm_1 <= MUX_v_32_2_2((line_buf3_Iy_rsci_q_d[31:0]),
          rdbuf3_Iy_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_31_itm_1 <= MUX_v_32_2_2((line_buf1_Iy_rsci_q_d[31:0]),
          rdbuf1_Iy_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_32_itm_1 <= MUX_v_32_2_2((line_buf0_Iy_rsci_q_d[31:0]),
          rdbuf0_Iy_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Iz0_lpi_1_dfm_1_2 <= Iz0_lpi_1_dfm_1_1;
      Gradient_weight_y_COLUMN_mux_33_itm_1 <= MUX_v_32_2_2((line_buf5_Iz_rsci_q_d[31:0]),
          rdbuf5_Iz_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_36_itm_1 <= MUX_v_32_2_2((line_buf2_Iz_rsci_q_d[31:0]),
          rdbuf2_Iz_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_34_itm_1 <= MUX_v_32_2_2((line_buf4_Iz_rsci_q_d[31:0]),
          rdbuf4_Iz_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_35_itm_1 <= MUX_v_32_2_2((line_buf3_Iz_rsci_q_d[31:0]),
          rdbuf3_Iz_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_37_itm_1 <= MUX_v_32_2_2((line_buf1_Iz_rsci_q_d[31:0]),
          rdbuf1_Iz_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_weight_y_COLUMN_mux_38_itm_1 <= MUX_v_32_2_2((line_buf0_Iz_rsci_q_d[31:0]),
          rdbuf0_Iz_lpi_1_63_32, Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      operator_9_false_1_slc_operator_9_false_1_acc_9_itm_1 <= readslicef_10_1_9(operator_9_false_1_acc_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      y_filtered_rsci_idat_95_64 <= 32'b00000000000000000000000000000000;
      y_filtered_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
      y_filtered_rsci_idat_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      y_filtered_rsci_idat_95_64 <= 32'b00000000000000000000000000000000;
      y_filtered_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
      y_filtered_rsci_idat_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( Gradient_weight_y_COLUMN_if_3_and_cse ) begin
      y_filtered_rsci_idat_95_64 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (readslicef_63_32_31(Gradient_weight_y_COLUMN_if_3_acc_21_nl)), Gradient_weight_y_COLUMN_if_3_not_3_nl);
      y_filtered_rsci_idat_31_0 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (readslicef_63_32_31(Gradient_weight_y_COLUMN_if_3_acc_nl)), Gradient_weight_y_COLUMN_if_3_not_4_nl);
      y_filtered_rsci_idat_63_32 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (readslicef_63_32_31(Gradient_weight_y_COLUMN_if_3_acc_20_nl)), Gradient_weight_y_COLUMN_if_3_not_5_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      wrbuf0_Iz_31_0_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      wrbuf0_Iy_31_0_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      wrbuf0_Ix_31_0_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      wrbuf0_Iz_31_0_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      wrbuf0_Iy_31_0_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      wrbuf0_Ix_31_0_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( wrbuf0_Iz_and_cse ) begin
      wrbuf0_Iz_31_0_lpi_1_dfm_2 <= wrbuf0_Iz_31_0_lpi_1_dfm_4;
      wrbuf0_Iy_31_0_lpi_1_dfm_2 <= wrbuf0_Iy_31_0_lpi_1_dfm_4;
      wrbuf0_Ix_31_0_lpi_1_dfm_2 <= wrbuf0_Ix_31_0_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rdbuf5_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf2_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf4_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf3_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf1_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf0_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf5_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf2_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf4_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf3_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf1_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf0_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf5_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf2_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf4_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf3_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf1_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf0_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      rdbuf5_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf2_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf4_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf3_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf1_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf0_Ix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf5_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf2_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf4_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf3_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf1_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf0_Iy_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf5_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf2_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf4_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf3_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf1_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf0_Iz_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( rdbuf5_Ix_and_cse ) begin
      rdbuf5_Ix_lpi_1_63_32 <= MUX_v_32_2_2(rdbuf5_Ix_lpi_1_dfm_1_63_32, (line_buf5_Ix_rsci_q_d[63:32]),
          and_dcpl_23);
      rdbuf2_Ix_lpi_1_63_32 <= MUX_v_32_2_2((line_buf2_Ix_rsci_q_d[63:32]), (rdbuf2_Ix_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf4_Ix_lpi_1_63_32 <= MUX_v_32_2_2((line_buf4_Ix_rsci_q_d[63:32]), (rdbuf4_Ix_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf3_Ix_lpi_1_63_32 <= MUX_v_32_2_2((line_buf3_Ix_rsci_q_d[63:32]), (rdbuf3_Ix_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf1_Ix_lpi_1_63_32 <= MUX_v_32_2_2((line_buf1_Ix_rsci_q_d[63:32]), (rdbuf1_Ix_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf0_Ix_lpi_1_63_32 <= MUX_v_32_2_2((line_buf0_Ix_rsci_q_d[63:32]), (rdbuf0_Ix_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf5_Iy_lpi_1_63_32 <= MUX_v_32_2_2(rdbuf5_Iy_lpi_1_dfm_1_63_32, (line_buf5_Iy_rsci_q_d[63:32]),
          and_dcpl_23);
      rdbuf2_Iy_lpi_1_63_32 <= MUX_v_32_2_2((line_buf2_Iy_rsci_q_d[63:32]), (rdbuf2_Iy_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf4_Iy_lpi_1_63_32 <= MUX_v_32_2_2((line_buf4_Iy_rsci_q_d[63:32]), (rdbuf4_Iy_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf3_Iy_lpi_1_63_32 <= MUX_v_32_2_2((line_buf3_Iy_rsci_q_d[63:32]), (rdbuf3_Iy_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf1_Iy_lpi_1_63_32 <= MUX_v_32_2_2((line_buf1_Iy_rsci_q_d[63:32]), (rdbuf1_Iy_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf0_Iy_lpi_1_63_32 <= MUX_v_32_2_2((line_buf0_Iy_rsci_q_d[63:32]), (rdbuf0_Iy_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf5_Iz_lpi_1_63_32 <= MUX_v_32_2_2(rdbuf5_Iz_lpi_1_dfm_1_63_32, (line_buf5_Iz_rsci_q_d[63:32]),
          and_dcpl_23);
      rdbuf2_Iz_lpi_1_63_32 <= MUX_v_32_2_2((line_buf2_Iz_rsci_q_d[63:32]), (rdbuf2_Iz_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf4_Iz_lpi_1_63_32 <= MUX_v_32_2_2((line_buf4_Iz_rsci_q_d[63:32]), (rdbuf4_Iz_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf3_Iz_lpi_1_63_32 <= MUX_v_32_2_2((line_buf3_Iz_rsci_q_d[63:32]), (rdbuf3_Iz_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf1_Iz_lpi_1_63_32 <= MUX_v_32_2_2((line_buf1_Iz_rsci_q_d[63:32]), (rdbuf1_Iz_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf0_Iz_lpi_1_63_32 <= MUX_v_32_2_2((line_buf0_Iz_rsci_q_d[63:32]), (rdbuf0_Iz_lpi_1_dfm_1[63:32]),
          Gradient_weight_y_COLUMN_x_lpi_1_dfm_2_0);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rdbuf5_Iz_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf5_Iy_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf5_Ix_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      rdbuf5_Iz_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf5_Iy_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf5_Ix_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( rdbuf5_Iz_and_1_cse ) begin
      rdbuf5_Iz_lpi_1_dfm_1_63_32 <= line_buf5_Iz_rsci_q_d[63:32];
      rdbuf5_Iy_lpi_1_dfm_1_63_32 <= line_buf5_Iy_rsci_q_d[63:32];
      rdbuf5_Ix_lpi_1_dfm_1_63_32 <= line_buf5_Ix_rsci_q_d[63:32];
    end
  end
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_27_itm_1  = conv_s2s_61_63(Gradient_weight_y_COLUMN_if_3_mul_15_itm_1)
      + conv_s2s_61_63({Gradient_weight_y_COLUMN_if_3_mul_16_itm_1 , 1'b0}) + conv_s2s_61_63({Gradient_weight_y_COLUMN_if_3_mul_18_itm_1
      , 1'b0}) + conv_s2s_61_63(Gradient_weight_y_COLUMN_if_3_mul_19_itm_1);
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_40_nl = (Gradient_weight_y_COLUMN_if_3_mul_20_itm_1[59:30])
      + 30'b000000000000000000000000000001;
  assign Gradient_weight_y_COLUMN_if_3_acc_40_nl = nl_Gradient_weight_y_COLUMN_if_3_acc_40_nl[29:0];
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_23_itm_1  = conv_s2s_60_61({Gradient_weight_y_COLUMN_if_3_acc_40_nl
      , (Gradient_weight_y_COLUMN_if_3_mul_20_itm_1[29:0])}) + conv_s2s_60_61(Gradient_weight_y_COLUMN_if_3_mul_14_itm_1);
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_39_itm_1  = conv_s2s_61_63(Gradient_weight_y_COLUMN_if_3_mul_1_itm_1)
      + conv_s2s_61_63({Gradient_weight_y_COLUMN_if_3_mul_2_itm_1 , 1'b0}) + conv_s2s_61_63({Gradient_weight_y_COLUMN_if_3_mul_4_itm_1
      , 1'b0}) + conv_s2s_61_63(Gradient_weight_y_COLUMN_if_3_mul_5_itm_1);
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_42_nl = (Gradient_weight_y_COLUMN_if_3_mul_6_itm_1[59:30])
      + 30'b000000000000000000000000000001;
  assign Gradient_weight_y_COLUMN_if_3_acc_42_nl = nl_Gradient_weight_y_COLUMN_if_3_acc_42_nl[29:0];
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_35_itm_1  = conv_s2s_60_61({Gradient_weight_y_COLUMN_if_3_acc_42_nl
      , (Gradient_weight_y_COLUMN_if_3_mul_6_itm_1[29:0])}) + conv_s2s_60_61(Gradient_weight_y_COLUMN_if_3_mul_itm_1);
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_33_itm_1  = conv_s2s_61_63(Gradient_weight_y_COLUMN_if_3_mul_8_itm_1)
      + conv_s2s_61_63({Gradient_weight_y_COLUMN_if_3_mul_9_itm_1 , 1'b0}) + conv_s2s_61_63({Gradient_weight_y_COLUMN_if_3_mul_11_itm_1
      , 1'b0}) + conv_s2s_61_63(Gradient_weight_y_COLUMN_if_3_mul_12_itm_1);
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_41_nl = (Gradient_weight_y_COLUMN_if_3_mul_13_itm_1[59:30])
      + 30'b000000000000000000000000000001;
  assign Gradient_weight_y_COLUMN_if_3_acc_41_nl = nl_Gradient_weight_y_COLUMN_if_3_acc_41_nl[29:0];
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_29_itm_1  = conv_s2s_60_61({Gradient_weight_y_COLUMN_if_3_acc_41_nl
      , (Gradient_weight_y_COLUMN_if_3_mul_13_itm_1[29:0])}) + conv_s2s_60_61(Gradient_weight_y_COLUMN_if_3_mul_7_itm_1);
  assign nl_Gradient_weight_y_COLUMN_aelse_acc_nl = ({1'b1 , Gradient_weight_y_ROW_y_lpi_1_dfm_2})
      + conv_u2u_9_10(~ heightIn) + 10'b0000000001;
  assign Gradient_weight_y_COLUMN_aelse_acc_nl = nl_Gradient_weight_y_COLUMN_aelse_acc_nl[9:0];
  assign nl_Gradient_weight_y_COLUMN_x_sva_2_1  = Gradient_weight_y_COLUMN_x_lpi_1_dfm_2
      + 11'b00000000001;
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_6_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_21_itm_1)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_itm_1  = $signed(Ix0_lpi_1_dfm_1_2)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_1_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_26_itm_1)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_2_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_25_itm_1)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_4_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_23_itm_1)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_5_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_22_itm_1)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_13_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_27_itm_1)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_7_itm_1  = $signed(Iy0_lpi_1_dfm_1_2)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_8_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_32_itm_1)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_9_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_31_itm_1)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_11_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_29_itm_1)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_12_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_28_itm_1)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_20_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_33_itm_1)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_14_itm_1  = $signed(Iz0_lpi_1_dfm_1_2)
      * $signed(29'b01001101010011111101111100111);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_15_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_38_itm_1)
      * $signed(30'b010001000001100010010011011101);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_16_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_37_itm_1)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_18_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_35_itm_1)
      * $signed(29'b01011111101100010101101101011);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_19_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_34_itm_1)
      * $signed(30'b010001000001100010010011011101);
  assign nl_operator_9_false_acc_nl = conv_u2u_8_9(Gradient_weight_y_ROW_y_lpi_1_dfm_1[8:1])
      + 9'b111111101;
  assign operator_9_false_acc_nl = nl_operator_9_false_acc_nl[8:0];
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_3_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_24_itm_1)
      * $signed(31'b0100101001010001000110011100111);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_10_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_30_itm_1)
      * $signed(31'b0100101001010001000110011100111);
  assign nl_Gradient_weight_y_COLUMN_if_3_mul_17_itm_1  = $signed(Gradient_weight_y_COLUMN_mux_36_itm_1)
      * $signed(31'b0100101001010001000110011100111);
  assign nl_operator_9_false_1_acc_nl = conv_u2s_9_10(Gradient_weight_y_ROW_y_lpi_1_dfm_2)
      + 10'b1111111101;
  assign operator_9_false_1_acc_nl = nl_operator_9_false_1_acc_nl[9:0];
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_26_nl = Gradient_weight_y_COLUMN_if_3_mul_17_itm_2
      + conv_s2s_61_62(Gradient_weight_y_COLUMN_if_3_acc_23_itm_1);
  assign Gradient_weight_y_COLUMN_if_3_acc_26_nl = nl_Gradient_weight_y_COLUMN_if_3_acc_26_nl[61:0];
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_21_nl = Gradient_weight_y_COLUMN_if_3_acc_27_itm_1
      + conv_s2s_62_63(Gradient_weight_y_COLUMN_if_3_acc_26_nl);
  assign Gradient_weight_y_COLUMN_if_3_acc_21_nl = nl_Gradient_weight_y_COLUMN_if_3_acc_21_nl[62:0];
  assign Gradient_weight_y_COLUMN_if_3_not_3_nl = ~ and_dcpl_21;
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_38_nl = Gradient_weight_y_COLUMN_if_3_mul_3_itm_2
      + conv_s2s_61_62(Gradient_weight_y_COLUMN_if_3_acc_35_itm_1);
  assign Gradient_weight_y_COLUMN_if_3_acc_38_nl = nl_Gradient_weight_y_COLUMN_if_3_acc_38_nl[61:0];
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_nl = Gradient_weight_y_COLUMN_if_3_acc_39_itm_1
      + conv_s2s_62_63(Gradient_weight_y_COLUMN_if_3_acc_38_nl);
  assign Gradient_weight_y_COLUMN_if_3_acc_nl = nl_Gradient_weight_y_COLUMN_if_3_acc_nl[62:0];
  assign Gradient_weight_y_COLUMN_if_3_not_4_nl = ~ and_dcpl_21;
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_32_nl = Gradient_weight_y_COLUMN_if_3_mul_10_itm_2
      + conv_s2s_61_62(Gradient_weight_y_COLUMN_if_3_acc_29_itm_1);
  assign Gradient_weight_y_COLUMN_if_3_acc_32_nl = nl_Gradient_weight_y_COLUMN_if_3_acc_32_nl[61:0];
  assign nl_Gradient_weight_y_COLUMN_if_3_acc_20_nl = Gradient_weight_y_COLUMN_if_3_acc_33_itm_1
      + conv_s2s_62_63(Gradient_weight_y_COLUMN_if_3_acc_32_nl);
  assign Gradient_weight_y_COLUMN_if_3_acc_20_nl = nl_Gradient_weight_y_COLUMN_if_3_acc_20_nl[62:0];
  assign Gradient_weight_y_COLUMN_if_3_not_5_nl = ~ and_dcpl_21;

  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [31:0] readslicef_63_32_31;
    input [62:0] vector;
    reg [62:0] tmp;
  begin
    tmp = vector >> 31;
    readslicef_63_32_31 = tmp[31:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [60:0] conv_s2s_60_61 ;
    input [59:0]  vector ;
  begin
    conv_s2s_60_61 = {vector[59], vector};
  end
  endfunction


  function automatic [61:0] conv_s2s_61_62 ;
    input [60:0]  vector ;
  begin
    conv_s2s_61_62 = {vector[60], vector};
  end
  endfunction


  function automatic [62:0] conv_s2s_61_63 ;
    input [60:0]  vector ;
  begin
    conv_s2s_61_63 = {{2{vector[60]}}, vector};
  end
  endfunction


  function automatic [62:0] conv_s2s_62_63 ;
    input [61:0]  vector ;
  begin
    conv_s2s_62_63 = {vector[61], vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y_struct
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y_struct (
  clk, rst, arst_n, gradient_x_rsc_dat, gradient_x_rsc_vld, gradient_x_rsc_rdy, gradient_y_rsc_dat,
      gradient_y_rsc_vld, gradient_y_rsc_rdy, gradient_z_rsc_dat, gradient_z_rsc_vld,
      gradient_z_rsc_rdy, y_filtered_rsc_dat_z, y_filtered_rsc_dat_y, y_filtered_rsc_dat_x,
      y_filtered_rsc_vld, y_filtered_rsc_rdy, widthIn, heightIn, line_buf5_Ix_rsc_clken,
      line_buf5_Ix_rsc_q, line_buf5_Ix_rsc_we, line_buf5_Ix_rsc_d, line_buf5_Ix_rsc_adr,
      line_buf4_Ix_rsc_clken, line_buf4_Ix_rsc_q, line_buf4_Ix_rsc_we, line_buf4_Ix_rsc_d,
      line_buf4_Ix_rsc_adr, line_buf3_Ix_rsc_clken, line_buf3_Ix_rsc_q, line_buf3_Ix_rsc_we,
      line_buf3_Ix_rsc_d, line_buf3_Ix_rsc_adr, line_buf2_Ix_rsc_clken, line_buf2_Ix_rsc_q,
      line_buf2_Ix_rsc_we, line_buf2_Ix_rsc_d, line_buf2_Ix_rsc_adr, line_buf1_Ix_rsc_clken,
      line_buf1_Ix_rsc_q, line_buf1_Ix_rsc_we, line_buf1_Ix_rsc_d, line_buf1_Ix_rsc_adr,
      line_buf0_Ix_rsc_clken, line_buf0_Ix_rsc_q, line_buf0_Ix_rsc_we, line_buf0_Ix_rsc_d,
      line_buf0_Ix_rsc_adr, line_buf5_Iy_rsc_clken, line_buf5_Iy_rsc_q, line_buf5_Iy_rsc_we,
      line_buf5_Iy_rsc_d, line_buf5_Iy_rsc_adr, line_buf4_Iy_rsc_clken, line_buf4_Iy_rsc_q,
      line_buf4_Iy_rsc_we, line_buf4_Iy_rsc_d, line_buf4_Iy_rsc_adr, line_buf3_Iy_rsc_clken,
      line_buf3_Iy_rsc_q, line_buf3_Iy_rsc_we, line_buf3_Iy_rsc_d, line_buf3_Iy_rsc_adr,
      line_buf2_Iy_rsc_clken, line_buf2_Iy_rsc_q, line_buf2_Iy_rsc_we, line_buf2_Iy_rsc_d,
      line_buf2_Iy_rsc_adr, line_buf1_Iy_rsc_clken, line_buf1_Iy_rsc_q, line_buf1_Iy_rsc_we,
      line_buf1_Iy_rsc_d, line_buf1_Iy_rsc_adr, line_buf0_Iy_rsc_clken, line_buf0_Iy_rsc_q,
      line_buf0_Iy_rsc_we, line_buf0_Iy_rsc_d, line_buf0_Iy_rsc_adr, line_buf5_Iz_rsc_clken,
      line_buf5_Iz_rsc_q, line_buf5_Iz_rsc_we, line_buf5_Iz_rsc_d, line_buf5_Iz_rsc_adr,
      line_buf4_Iz_rsc_clken, line_buf4_Iz_rsc_q, line_buf4_Iz_rsc_we, line_buf4_Iz_rsc_d,
      line_buf4_Iz_rsc_adr, line_buf3_Iz_rsc_clken, line_buf3_Iz_rsc_q, line_buf3_Iz_rsc_we,
      line_buf3_Iz_rsc_d, line_buf3_Iz_rsc_adr, line_buf2_Iz_rsc_clken, line_buf2_Iz_rsc_q,
      line_buf2_Iz_rsc_we, line_buf2_Iz_rsc_d, line_buf2_Iz_rsc_adr, line_buf1_Iz_rsc_clken,
      line_buf1_Iz_rsc_q, line_buf1_Iz_rsc_we, line_buf1_Iz_rsc_d, line_buf1_Iz_rsc_adr,
      line_buf0_Iz_rsc_clken, line_buf0_Iz_rsc_q, line_buf0_Iz_rsc_we, line_buf0_Iz_rsc_d,
      line_buf0_Iz_rsc_adr
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] gradient_x_rsc_dat;
  input gradient_x_rsc_vld;
  output gradient_x_rsc_rdy;
  input [31:0] gradient_y_rsc_dat;
  input gradient_y_rsc_vld;
  output gradient_y_rsc_rdy;
  input [31:0] gradient_z_rsc_dat;
  input gradient_z_rsc_vld;
  output gradient_z_rsc_rdy;
  output [31:0] y_filtered_rsc_dat_z;
  output [31:0] y_filtered_rsc_dat_y;
  output [31:0] y_filtered_rsc_dat_x;
  output y_filtered_rsc_vld;
  input y_filtered_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  output line_buf5_Ix_rsc_clken;
  input [63:0] line_buf5_Ix_rsc_q;
  output line_buf5_Ix_rsc_we;
  output [63:0] line_buf5_Ix_rsc_d;
  output [8:0] line_buf5_Ix_rsc_adr;
  output line_buf4_Ix_rsc_clken;
  input [63:0] line_buf4_Ix_rsc_q;
  output line_buf4_Ix_rsc_we;
  output [63:0] line_buf4_Ix_rsc_d;
  output [8:0] line_buf4_Ix_rsc_adr;
  output line_buf3_Ix_rsc_clken;
  input [63:0] line_buf3_Ix_rsc_q;
  output line_buf3_Ix_rsc_we;
  output [63:0] line_buf3_Ix_rsc_d;
  output [8:0] line_buf3_Ix_rsc_adr;
  output line_buf2_Ix_rsc_clken;
  input [63:0] line_buf2_Ix_rsc_q;
  output line_buf2_Ix_rsc_we;
  output [63:0] line_buf2_Ix_rsc_d;
  output [8:0] line_buf2_Ix_rsc_adr;
  output line_buf1_Ix_rsc_clken;
  input [63:0] line_buf1_Ix_rsc_q;
  output line_buf1_Ix_rsc_we;
  output [63:0] line_buf1_Ix_rsc_d;
  output [8:0] line_buf1_Ix_rsc_adr;
  output line_buf0_Ix_rsc_clken;
  input [63:0] line_buf0_Ix_rsc_q;
  output line_buf0_Ix_rsc_we;
  output [63:0] line_buf0_Ix_rsc_d;
  output [8:0] line_buf0_Ix_rsc_adr;
  output line_buf5_Iy_rsc_clken;
  input [63:0] line_buf5_Iy_rsc_q;
  output line_buf5_Iy_rsc_we;
  output [63:0] line_buf5_Iy_rsc_d;
  output [8:0] line_buf5_Iy_rsc_adr;
  output line_buf4_Iy_rsc_clken;
  input [63:0] line_buf4_Iy_rsc_q;
  output line_buf4_Iy_rsc_we;
  output [63:0] line_buf4_Iy_rsc_d;
  output [8:0] line_buf4_Iy_rsc_adr;
  output line_buf3_Iy_rsc_clken;
  input [63:0] line_buf3_Iy_rsc_q;
  output line_buf3_Iy_rsc_we;
  output [63:0] line_buf3_Iy_rsc_d;
  output [8:0] line_buf3_Iy_rsc_adr;
  output line_buf2_Iy_rsc_clken;
  input [63:0] line_buf2_Iy_rsc_q;
  output line_buf2_Iy_rsc_we;
  output [63:0] line_buf2_Iy_rsc_d;
  output [8:0] line_buf2_Iy_rsc_adr;
  output line_buf1_Iy_rsc_clken;
  input [63:0] line_buf1_Iy_rsc_q;
  output line_buf1_Iy_rsc_we;
  output [63:0] line_buf1_Iy_rsc_d;
  output [8:0] line_buf1_Iy_rsc_adr;
  output line_buf0_Iy_rsc_clken;
  input [63:0] line_buf0_Iy_rsc_q;
  output line_buf0_Iy_rsc_we;
  output [63:0] line_buf0_Iy_rsc_d;
  output [8:0] line_buf0_Iy_rsc_adr;
  output line_buf5_Iz_rsc_clken;
  input [63:0] line_buf5_Iz_rsc_q;
  output line_buf5_Iz_rsc_we;
  output [63:0] line_buf5_Iz_rsc_d;
  output [8:0] line_buf5_Iz_rsc_adr;
  output line_buf4_Iz_rsc_clken;
  input [63:0] line_buf4_Iz_rsc_q;
  output line_buf4_Iz_rsc_we;
  output [63:0] line_buf4_Iz_rsc_d;
  output [8:0] line_buf4_Iz_rsc_adr;
  output line_buf3_Iz_rsc_clken;
  input [63:0] line_buf3_Iz_rsc_q;
  output line_buf3_Iz_rsc_we;
  output [63:0] line_buf3_Iz_rsc_d;
  output [8:0] line_buf3_Iz_rsc_adr;
  output line_buf2_Iz_rsc_clken;
  input [63:0] line_buf2_Iz_rsc_q;
  output line_buf2_Iz_rsc_we;
  output [63:0] line_buf2_Iz_rsc_d;
  output [8:0] line_buf2_Iz_rsc_adr;
  output line_buf1_Iz_rsc_clken;
  input [63:0] line_buf1_Iz_rsc_q;
  output line_buf1_Iz_rsc_we;
  output [63:0] line_buf1_Iz_rsc_d;
  output [8:0] line_buf1_Iz_rsc_adr;
  output line_buf0_Iz_rsc_clken;
  input [63:0] line_buf0_Iz_rsc_q;
  output line_buf0_Iz_rsc_we;
  output [63:0] line_buf0_Iz_rsc_d;
  output [8:0] line_buf0_Iz_rsc_adr;


  // Interconnect Declarations
  wire line_buf5_Ix_rsci_clken_d;
  wire [63:0] line_buf5_Ix_rsci_d_d;
  wire [63:0] line_buf5_Ix_rsci_q_d;
  wire [63:0] line_buf4_Ix_rsci_d_d;
  wire [63:0] line_buf4_Ix_rsci_q_d;
  wire [63:0] line_buf3_Ix_rsci_d_d;
  wire [63:0] line_buf3_Ix_rsci_q_d;
  wire [63:0] line_buf2_Ix_rsci_d_d;
  wire [63:0] line_buf2_Ix_rsci_q_d;
  wire [63:0] line_buf1_Ix_rsci_d_d;
  wire [63:0] line_buf1_Ix_rsci_q_d;
  wire [63:0] line_buf0_Ix_rsci_d_d;
  wire [63:0] line_buf0_Ix_rsci_q_d;
  wire [63:0] line_buf5_Iy_rsci_d_d;
  wire [63:0] line_buf5_Iy_rsci_q_d;
  wire [63:0] line_buf4_Iy_rsci_d_d;
  wire [63:0] line_buf4_Iy_rsci_q_d;
  wire [63:0] line_buf3_Iy_rsci_d_d;
  wire [63:0] line_buf3_Iy_rsci_q_d;
  wire [63:0] line_buf2_Iy_rsci_d_d;
  wire [63:0] line_buf2_Iy_rsci_q_d;
  wire [63:0] line_buf1_Iy_rsci_d_d;
  wire [63:0] line_buf1_Iy_rsci_q_d;
  wire [63:0] line_buf0_Iy_rsci_d_d;
  wire [63:0] line_buf0_Iy_rsci_q_d;
  wire [63:0] line_buf5_Iz_rsci_d_d;
  wire [63:0] line_buf5_Iz_rsci_q_d;
  wire [63:0] line_buf4_Iz_rsci_d_d;
  wire [63:0] line_buf4_Iz_rsci_q_d;
  wire [63:0] line_buf3_Iz_rsci_d_d;
  wire [63:0] line_buf3_Iz_rsci_q_d;
  wire [63:0] line_buf2_Iz_rsci_d_d;
  wire [63:0] line_buf2_Iz_rsci_q_d;
  wire [63:0] line_buf1_Iz_rsci_d_d;
  wire [63:0] line_buf1_Iz_rsci_q_d;
  wire [63:0] line_buf0_Iz_rsci_d_d;
  wire [63:0] line_buf0_Iz_rsci_q_d;
  wire [95:0] y_filtered_rsc_dat;
  wire [8:0] line_buf5_Ix_rsci_adr_d_iff;
  wire line_buf5_Ix_rsci_we_d_iff;
  wire line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff;


  // Interconnect Declarations for Component Instantiations 
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_7_9_64_512_1_512_64_1_gen
      line_buf5_Ix_rsci (
      .clken(line_buf5_Ix_rsc_clken),
      .q(line_buf5_Ix_rsc_q),
      .we(line_buf5_Ix_rsc_we),
      .d(line_buf5_Ix_rsc_d),
      .adr(line_buf5_Ix_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf5_Ix_rsci_d_d),
      .q_d(line_buf5_Ix_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_8_9_64_512_1_512_64_1_gen
      line_buf4_Ix_rsci (
      .clken(line_buf4_Ix_rsc_clken),
      .q(line_buf4_Ix_rsc_q),
      .we(line_buf4_Ix_rsc_we),
      .d(line_buf4_Ix_rsc_d),
      .adr(line_buf4_Ix_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf4_Ix_rsci_d_d),
      .q_d(line_buf4_Ix_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_9_9_64_512_1_512_64_1_gen
      line_buf3_Ix_rsci (
      .clken(line_buf3_Ix_rsc_clken),
      .q(line_buf3_Ix_rsc_q),
      .we(line_buf3_Ix_rsc_we),
      .d(line_buf3_Ix_rsc_d),
      .adr(line_buf3_Ix_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf3_Ix_rsci_d_d),
      .q_d(line_buf3_Ix_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_10_9_64_512_1_512_64_1_gen
      line_buf2_Ix_rsci (
      .clken(line_buf2_Ix_rsc_clken),
      .q(line_buf2_Ix_rsc_q),
      .we(line_buf2_Ix_rsc_we),
      .d(line_buf2_Ix_rsc_d),
      .adr(line_buf2_Ix_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf2_Ix_rsci_d_d),
      .q_d(line_buf2_Ix_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_11_9_64_512_1_512_64_1_gen
      line_buf1_Ix_rsci (
      .clken(line_buf1_Ix_rsc_clken),
      .q(line_buf1_Ix_rsc_q),
      .we(line_buf1_Ix_rsc_we),
      .d(line_buf1_Ix_rsc_d),
      .adr(line_buf1_Ix_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf1_Ix_rsci_d_d),
      .q_d(line_buf1_Ix_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_12_9_64_512_1_512_64_1_gen
      line_buf0_Ix_rsci (
      .clken(line_buf0_Ix_rsc_clken),
      .q(line_buf0_Ix_rsc_q),
      .we(line_buf0_Ix_rsc_we),
      .d(line_buf0_Ix_rsc_d),
      .adr(line_buf0_Ix_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf0_Ix_rsci_d_d),
      .q_d(line_buf0_Ix_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_13_9_64_512_1_512_64_1_gen
      line_buf5_Iy_rsci (
      .clken(line_buf5_Iy_rsc_clken),
      .q(line_buf5_Iy_rsc_q),
      .we(line_buf5_Iy_rsc_we),
      .d(line_buf5_Iy_rsc_d),
      .adr(line_buf5_Iy_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf5_Iy_rsci_d_d),
      .q_d(line_buf5_Iy_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_14_9_64_512_1_512_64_1_gen
      line_buf4_Iy_rsci (
      .clken(line_buf4_Iy_rsc_clken),
      .q(line_buf4_Iy_rsc_q),
      .we(line_buf4_Iy_rsc_we),
      .d(line_buf4_Iy_rsc_d),
      .adr(line_buf4_Iy_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf4_Iy_rsci_d_d),
      .q_d(line_buf4_Iy_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_15_9_64_512_1_512_64_1_gen
      line_buf3_Iy_rsci (
      .clken(line_buf3_Iy_rsc_clken),
      .q(line_buf3_Iy_rsc_q),
      .we(line_buf3_Iy_rsc_we),
      .d(line_buf3_Iy_rsc_d),
      .adr(line_buf3_Iy_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf3_Iy_rsci_d_d),
      .q_d(line_buf3_Iy_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_16_9_64_512_1_512_64_1_gen
      line_buf2_Iy_rsci (
      .clken(line_buf2_Iy_rsc_clken),
      .q(line_buf2_Iy_rsc_q),
      .we(line_buf2_Iy_rsc_we),
      .d(line_buf2_Iy_rsc_d),
      .adr(line_buf2_Iy_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf2_Iy_rsci_d_d),
      .q_d(line_buf2_Iy_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_17_9_64_512_1_512_64_1_gen
      line_buf1_Iy_rsci (
      .clken(line_buf1_Iy_rsc_clken),
      .q(line_buf1_Iy_rsc_q),
      .we(line_buf1_Iy_rsc_we),
      .d(line_buf1_Iy_rsc_d),
      .adr(line_buf1_Iy_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf1_Iy_rsci_d_d),
      .q_d(line_buf1_Iy_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_18_9_64_512_1_512_64_1_gen
      line_buf0_Iy_rsci (
      .clken(line_buf0_Iy_rsc_clken),
      .q(line_buf0_Iy_rsc_q),
      .we(line_buf0_Iy_rsc_we),
      .d(line_buf0_Iy_rsc_d),
      .adr(line_buf0_Iy_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf0_Iy_rsci_d_d),
      .q_d(line_buf0_Iy_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_19_9_64_512_1_512_64_1_gen
      line_buf5_Iz_rsci (
      .clken(line_buf5_Iz_rsc_clken),
      .q(line_buf5_Iz_rsc_q),
      .we(line_buf5_Iz_rsc_we),
      .d(line_buf5_Iz_rsc_d),
      .adr(line_buf5_Iz_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf5_Iz_rsci_d_d),
      .q_d(line_buf5_Iz_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_20_9_64_512_1_512_64_1_gen
      line_buf4_Iz_rsci (
      .clken(line_buf4_Iz_rsc_clken),
      .q(line_buf4_Iz_rsc_q),
      .we(line_buf4_Iz_rsc_we),
      .d(line_buf4_Iz_rsc_d),
      .adr(line_buf4_Iz_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf4_Iz_rsci_d_d),
      .q_d(line_buf4_Iz_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_21_9_64_512_1_512_64_1_gen
      line_buf3_Iz_rsci (
      .clken(line_buf3_Iz_rsc_clken),
      .q(line_buf3_Iz_rsc_q),
      .we(line_buf3_Iz_rsc_we),
      .d(line_buf3_Iz_rsc_d),
      .adr(line_buf3_Iz_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf3_Iz_rsci_d_d),
      .q_d(line_buf3_Iz_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_22_9_64_512_1_512_64_1_gen
      line_buf2_Iz_rsci (
      .clken(line_buf2_Iz_rsc_clken),
      .q(line_buf2_Iz_rsc_q),
      .we(line_buf2_Iz_rsc_we),
      .d(line_buf2_Iz_rsc_d),
      .adr(line_buf2_Iz_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf2_Iz_rsci_d_d),
      .q_d(line_buf2_Iz_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_23_9_64_512_1_512_64_1_gen
      line_buf1_Iz_rsci (
      .clken(line_buf1_Iz_rsc_clken),
      .q(line_buf1_Iz_rsc_q),
      .we(line_buf1_Iz_rsc_we),
      .d(line_buf1_Iz_rsc_d),
      .adr(line_buf1_Iz_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf1_Iz_rsci_d_d),
      .q_d(line_buf1_Iz_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_24_9_64_512_1_512_64_1_gen
      line_buf0_Iz_rsci (
      .clken(line_buf0_Iz_rsc_clken),
      .q(line_buf0_Iz_rsc_q),
      .we(line_buf0_Iz_rsc_we),
      .d(line_buf0_Iz_rsc_d),
      .adr(line_buf0_Iz_rsc_adr),
      .adr_d(line_buf5_Ix_rsci_adr_d_iff),
      .clken_d(line_buf5_Ix_rsci_clken_d),
      .d_d(line_buf0_Iz_rsci_d_d),
      .q_d(line_buf0_Iz_rsci_q_d),
      .we_d(line_buf5_Ix_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf5_Ix_rsci_we_d_iff)
    );
  OpticalFlow_gradient_weight_y_run OpticalFlow_gradient_weight_y_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .gradient_x_rsc_dat(gradient_x_rsc_dat),
      .gradient_x_rsc_vld(gradient_x_rsc_vld),
      .gradient_x_rsc_rdy(gradient_x_rsc_rdy),
      .gradient_y_rsc_dat(gradient_y_rsc_dat),
      .gradient_y_rsc_vld(gradient_y_rsc_vld),
      .gradient_y_rsc_rdy(gradient_y_rsc_rdy),
      .gradient_z_rsc_dat(gradient_z_rsc_dat),
      .gradient_z_rsc_vld(gradient_z_rsc_vld),
      .gradient_z_rsc_rdy(gradient_z_rsc_rdy),
      .y_filtered_rsc_dat(y_filtered_rsc_dat),
      .y_filtered_rsc_vld(y_filtered_rsc_vld),
      .y_filtered_rsc_rdy(y_filtered_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .line_buf5_Ix_rsci_clken_d(line_buf5_Ix_rsci_clken_d),
      .line_buf5_Ix_rsci_d_d(line_buf5_Ix_rsci_d_d),
      .line_buf5_Ix_rsci_q_d(line_buf5_Ix_rsci_q_d),
      .line_buf4_Ix_rsci_d_d(line_buf4_Ix_rsci_d_d),
      .line_buf4_Ix_rsci_q_d(line_buf4_Ix_rsci_q_d),
      .line_buf3_Ix_rsci_d_d(line_buf3_Ix_rsci_d_d),
      .line_buf3_Ix_rsci_q_d(line_buf3_Ix_rsci_q_d),
      .line_buf2_Ix_rsci_d_d(line_buf2_Ix_rsci_d_d),
      .line_buf2_Ix_rsci_q_d(line_buf2_Ix_rsci_q_d),
      .line_buf1_Ix_rsci_d_d(line_buf1_Ix_rsci_d_d),
      .line_buf1_Ix_rsci_q_d(line_buf1_Ix_rsci_q_d),
      .line_buf0_Ix_rsci_d_d(line_buf0_Ix_rsci_d_d),
      .line_buf0_Ix_rsci_q_d(line_buf0_Ix_rsci_q_d),
      .line_buf5_Iy_rsci_d_d(line_buf5_Iy_rsci_d_d),
      .line_buf5_Iy_rsci_q_d(line_buf5_Iy_rsci_q_d),
      .line_buf4_Iy_rsci_d_d(line_buf4_Iy_rsci_d_d),
      .line_buf4_Iy_rsci_q_d(line_buf4_Iy_rsci_q_d),
      .line_buf3_Iy_rsci_d_d(line_buf3_Iy_rsci_d_d),
      .line_buf3_Iy_rsci_q_d(line_buf3_Iy_rsci_q_d),
      .line_buf2_Iy_rsci_d_d(line_buf2_Iy_rsci_d_d),
      .line_buf2_Iy_rsci_q_d(line_buf2_Iy_rsci_q_d),
      .line_buf1_Iy_rsci_d_d(line_buf1_Iy_rsci_d_d),
      .line_buf1_Iy_rsci_q_d(line_buf1_Iy_rsci_q_d),
      .line_buf0_Iy_rsci_d_d(line_buf0_Iy_rsci_d_d),
      .line_buf0_Iy_rsci_q_d(line_buf0_Iy_rsci_q_d),
      .line_buf5_Iz_rsci_d_d(line_buf5_Iz_rsci_d_d),
      .line_buf5_Iz_rsci_q_d(line_buf5_Iz_rsci_q_d),
      .line_buf4_Iz_rsci_d_d(line_buf4_Iz_rsci_d_d),
      .line_buf4_Iz_rsci_q_d(line_buf4_Iz_rsci_q_d),
      .line_buf3_Iz_rsci_d_d(line_buf3_Iz_rsci_d_d),
      .line_buf3_Iz_rsci_q_d(line_buf3_Iz_rsci_q_d),
      .line_buf2_Iz_rsci_d_d(line_buf2_Iz_rsci_d_d),
      .line_buf2_Iz_rsci_q_d(line_buf2_Iz_rsci_q_d),
      .line_buf1_Iz_rsci_d_d(line_buf1_Iz_rsci_d_d),
      .line_buf1_Iz_rsci_q_d(line_buf1_Iz_rsci_q_d),
      .line_buf0_Iz_rsci_d_d(line_buf0_Iz_rsci_d_d),
      .line_buf0_Iz_rsci_q_d(line_buf0_Iz_rsci_q_d),
      .line_buf5_Ix_rsci_adr_d_pff(line_buf5_Ix_rsci_adr_d_iff),
      .line_buf5_Ix_rsci_we_d_pff(line_buf5_Ix_rsci_we_d_iff),
      .line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff(line_buf5_Ix_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff)
    );
  assign y_filtered_rsc_dat_x = y_filtered_rsc_dat[31:0];
  assign y_filtered_rsc_dat_y = y_filtered_rsc_dat[63:32];
  assign y_filtered_rsc_dat_z = y_filtered_rsc_dat[95:64];
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_weight_y
// ------------------------------------------------------------------


module OpticalFlow_gradient_weight_y (
  clk, rst, arst_n, gradient_x_rsc_dat, gradient_x_rsc_vld, gradient_x_rsc_rdy, gradient_y_rsc_dat,
      gradient_y_rsc_vld, gradient_y_rsc_rdy, gradient_z_rsc_dat, gradient_z_rsc_vld,
      gradient_z_rsc_rdy, y_filtered_rsc_dat, y_filtered_rsc_vld, y_filtered_rsc_rdy,
      widthIn, heightIn, line_buf5_Ix_rsc_clken, line_buf5_Ix_rsc_q, line_buf5_Ix_rsc_we,
      line_buf5_Ix_rsc_d, line_buf5_Ix_rsc_adr, line_buf4_Ix_rsc_clken, line_buf4_Ix_rsc_q,
      line_buf4_Ix_rsc_we, line_buf4_Ix_rsc_d, line_buf4_Ix_rsc_adr, line_buf3_Ix_rsc_clken,
      line_buf3_Ix_rsc_q, line_buf3_Ix_rsc_we, line_buf3_Ix_rsc_d, line_buf3_Ix_rsc_adr,
      line_buf2_Ix_rsc_clken, line_buf2_Ix_rsc_q, line_buf2_Ix_rsc_we, line_buf2_Ix_rsc_d,
      line_buf2_Ix_rsc_adr, line_buf1_Ix_rsc_clken, line_buf1_Ix_rsc_q, line_buf1_Ix_rsc_we,
      line_buf1_Ix_rsc_d, line_buf1_Ix_rsc_adr, line_buf0_Ix_rsc_clken, line_buf0_Ix_rsc_q,
      line_buf0_Ix_rsc_we, line_buf0_Ix_rsc_d, line_buf0_Ix_rsc_adr, line_buf5_Iy_rsc_clken,
      line_buf5_Iy_rsc_q, line_buf5_Iy_rsc_we, line_buf5_Iy_rsc_d, line_buf5_Iy_rsc_adr,
      line_buf4_Iy_rsc_clken, line_buf4_Iy_rsc_q, line_buf4_Iy_rsc_we, line_buf4_Iy_rsc_d,
      line_buf4_Iy_rsc_adr, line_buf3_Iy_rsc_clken, line_buf3_Iy_rsc_q, line_buf3_Iy_rsc_we,
      line_buf3_Iy_rsc_d, line_buf3_Iy_rsc_adr, line_buf2_Iy_rsc_clken, line_buf2_Iy_rsc_q,
      line_buf2_Iy_rsc_we, line_buf2_Iy_rsc_d, line_buf2_Iy_rsc_adr, line_buf1_Iy_rsc_clken,
      line_buf1_Iy_rsc_q, line_buf1_Iy_rsc_we, line_buf1_Iy_rsc_d, line_buf1_Iy_rsc_adr,
      line_buf0_Iy_rsc_clken, line_buf0_Iy_rsc_q, line_buf0_Iy_rsc_we, line_buf0_Iy_rsc_d,
      line_buf0_Iy_rsc_adr, line_buf5_Iz_rsc_clken, line_buf5_Iz_rsc_q, line_buf5_Iz_rsc_we,
      line_buf5_Iz_rsc_d, line_buf5_Iz_rsc_adr, line_buf4_Iz_rsc_clken, line_buf4_Iz_rsc_q,
      line_buf4_Iz_rsc_we, line_buf4_Iz_rsc_d, line_buf4_Iz_rsc_adr, line_buf3_Iz_rsc_clken,
      line_buf3_Iz_rsc_q, line_buf3_Iz_rsc_we, line_buf3_Iz_rsc_d, line_buf3_Iz_rsc_adr,
      line_buf2_Iz_rsc_clken, line_buf2_Iz_rsc_q, line_buf2_Iz_rsc_we, line_buf2_Iz_rsc_d,
      line_buf2_Iz_rsc_adr, line_buf1_Iz_rsc_clken, line_buf1_Iz_rsc_q, line_buf1_Iz_rsc_we,
      line_buf1_Iz_rsc_d, line_buf1_Iz_rsc_adr, line_buf0_Iz_rsc_clken, line_buf0_Iz_rsc_q,
      line_buf0_Iz_rsc_we, line_buf0_Iz_rsc_d, line_buf0_Iz_rsc_adr
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] gradient_x_rsc_dat;
  input gradient_x_rsc_vld;
  output gradient_x_rsc_rdy;
  input [31:0] gradient_y_rsc_dat;
  input gradient_y_rsc_vld;
  output gradient_y_rsc_rdy;
  input [31:0] gradient_z_rsc_dat;
  input gradient_z_rsc_vld;
  output gradient_z_rsc_rdy;
  output [95:0] y_filtered_rsc_dat;
  output y_filtered_rsc_vld;
  input y_filtered_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  output line_buf5_Ix_rsc_clken;
  input [63:0] line_buf5_Ix_rsc_q;
  output line_buf5_Ix_rsc_we;
  output [63:0] line_buf5_Ix_rsc_d;
  output [8:0] line_buf5_Ix_rsc_adr;
  output line_buf4_Ix_rsc_clken;
  input [63:0] line_buf4_Ix_rsc_q;
  output line_buf4_Ix_rsc_we;
  output [63:0] line_buf4_Ix_rsc_d;
  output [8:0] line_buf4_Ix_rsc_adr;
  output line_buf3_Ix_rsc_clken;
  input [63:0] line_buf3_Ix_rsc_q;
  output line_buf3_Ix_rsc_we;
  output [63:0] line_buf3_Ix_rsc_d;
  output [8:0] line_buf3_Ix_rsc_adr;
  output line_buf2_Ix_rsc_clken;
  input [63:0] line_buf2_Ix_rsc_q;
  output line_buf2_Ix_rsc_we;
  output [63:0] line_buf2_Ix_rsc_d;
  output [8:0] line_buf2_Ix_rsc_adr;
  output line_buf1_Ix_rsc_clken;
  input [63:0] line_buf1_Ix_rsc_q;
  output line_buf1_Ix_rsc_we;
  output [63:0] line_buf1_Ix_rsc_d;
  output [8:0] line_buf1_Ix_rsc_adr;
  output line_buf0_Ix_rsc_clken;
  input [63:0] line_buf0_Ix_rsc_q;
  output line_buf0_Ix_rsc_we;
  output [63:0] line_buf0_Ix_rsc_d;
  output [8:0] line_buf0_Ix_rsc_adr;
  output line_buf5_Iy_rsc_clken;
  input [63:0] line_buf5_Iy_rsc_q;
  output line_buf5_Iy_rsc_we;
  output [63:0] line_buf5_Iy_rsc_d;
  output [8:0] line_buf5_Iy_rsc_adr;
  output line_buf4_Iy_rsc_clken;
  input [63:0] line_buf4_Iy_rsc_q;
  output line_buf4_Iy_rsc_we;
  output [63:0] line_buf4_Iy_rsc_d;
  output [8:0] line_buf4_Iy_rsc_adr;
  output line_buf3_Iy_rsc_clken;
  input [63:0] line_buf3_Iy_rsc_q;
  output line_buf3_Iy_rsc_we;
  output [63:0] line_buf3_Iy_rsc_d;
  output [8:0] line_buf3_Iy_rsc_adr;
  output line_buf2_Iy_rsc_clken;
  input [63:0] line_buf2_Iy_rsc_q;
  output line_buf2_Iy_rsc_we;
  output [63:0] line_buf2_Iy_rsc_d;
  output [8:0] line_buf2_Iy_rsc_adr;
  output line_buf1_Iy_rsc_clken;
  input [63:0] line_buf1_Iy_rsc_q;
  output line_buf1_Iy_rsc_we;
  output [63:0] line_buf1_Iy_rsc_d;
  output [8:0] line_buf1_Iy_rsc_adr;
  output line_buf0_Iy_rsc_clken;
  input [63:0] line_buf0_Iy_rsc_q;
  output line_buf0_Iy_rsc_we;
  output [63:0] line_buf0_Iy_rsc_d;
  output [8:0] line_buf0_Iy_rsc_adr;
  output line_buf5_Iz_rsc_clken;
  input [63:0] line_buf5_Iz_rsc_q;
  output line_buf5_Iz_rsc_we;
  output [63:0] line_buf5_Iz_rsc_d;
  output [8:0] line_buf5_Iz_rsc_adr;
  output line_buf4_Iz_rsc_clken;
  input [63:0] line_buf4_Iz_rsc_q;
  output line_buf4_Iz_rsc_we;
  output [63:0] line_buf4_Iz_rsc_d;
  output [8:0] line_buf4_Iz_rsc_adr;
  output line_buf3_Iz_rsc_clken;
  input [63:0] line_buf3_Iz_rsc_q;
  output line_buf3_Iz_rsc_we;
  output [63:0] line_buf3_Iz_rsc_d;
  output [8:0] line_buf3_Iz_rsc_adr;
  output line_buf2_Iz_rsc_clken;
  input [63:0] line_buf2_Iz_rsc_q;
  output line_buf2_Iz_rsc_we;
  output [63:0] line_buf2_Iz_rsc_d;
  output [8:0] line_buf2_Iz_rsc_adr;
  output line_buf1_Iz_rsc_clken;
  input [63:0] line_buf1_Iz_rsc_q;
  output line_buf1_Iz_rsc_we;
  output [63:0] line_buf1_Iz_rsc_d;
  output [8:0] line_buf1_Iz_rsc_adr;
  output line_buf0_Iz_rsc_clken;
  input [63:0] line_buf0_Iz_rsc_q;
  output line_buf0_Iz_rsc_we;
  output [63:0] line_buf0_Iz_rsc_d;
  output [8:0] line_buf0_Iz_rsc_adr;


  // Interconnect Declarations
  wire [31:0] y_filtered_rsc_dat_z;
  wire [31:0] y_filtered_rsc_dat_y;
  wire [31:0] y_filtered_rsc_dat_x;


  // Interconnect Declarations for Component Instantiations 
  OpticalFlow_gradient_weight_y_struct OpticalFlow_gradient_weight_y_struct_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .gradient_x_rsc_dat(gradient_x_rsc_dat),
      .gradient_x_rsc_vld(gradient_x_rsc_vld),
      .gradient_x_rsc_rdy(gradient_x_rsc_rdy),
      .gradient_y_rsc_dat(gradient_y_rsc_dat),
      .gradient_y_rsc_vld(gradient_y_rsc_vld),
      .gradient_y_rsc_rdy(gradient_y_rsc_rdy),
      .gradient_z_rsc_dat(gradient_z_rsc_dat),
      .gradient_z_rsc_vld(gradient_z_rsc_vld),
      .gradient_z_rsc_rdy(gradient_z_rsc_rdy),
      .y_filtered_rsc_dat_z(y_filtered_rsc_dat_z),
      .y_filtered_rsc_dat_y(y_filtered_rsc_dat_y),
      .y_filtered_rsc_dat_x(y_filtered_rsc_dat_x),
      .y_filtered_rsc_vld(y_filtered_rsc_vld),
      .y_filtered_rsc_rdy(y_filtered_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .line_buf5_Ix_rsc_clken(line_buf5_Ix_rsc_clken),
      .line_buf5_Ix_rsc_q(line_buf5_Ix_rsc_q),
      .line_buf5_Ix_rsc_we(line_buf5_Ix_rsc_we),
      .line_buf5_Ix_rsc_d(line_buf5_Ix_rsc_d),
      .line_buf5_Ix_rsc_adr(line_buf5_Ix_rsc_adr),
      .line_buf4_Ix_rsc_clken(line_buf4_Ix_rsc_clken),
      .line_buf4_Ix_rsc_q(line_buf4_Ix_rsc_q),
      .line_buf4_Ix_rsc_we(line_buf4_Ix_rsc_we),
      .line_buf4_Ix_rsc_d(line_buf4_Ix_rsc_d),
      .line_buf4_Ix_rsc_adr(line_buf4_Ix_rsc_adr),
      .line_buf3_Ix_rsc_clken(line_buf3_Ix_rsc_clken),
      .line_buf3_Ix_rsc_q(line_buf3_Ix_rsc_q),
      .line_buf3_Ix_rsc_we(line_buf3_Ix_rsc_we),
      .line_buf3_Ix_rsc_d(line_buf3_Ix_rsc_d),
      .line_buf3_Ix_rsc_adr(line_buf3_Ix_rsc_adr),
      .line_buf2_Ix_rsc_clken(line_buf2_Ix_rsc_clken),
      .line_buf2_Ix_rsc_q(line_buf2_Ix_rsc_q),
      .line_buf2_Ix_rsc_we(line_buf2_Ix_rsc_we),
      .line_buf2_Ix_rsc_d(line_buf2_Ix_rsc_d),
      .line_buf2_Ix_rsc_adr(line_buf2_Ix_rsc_adr),
      .line_buf1_Ix_rsc_clken(line_buf1_Ix_rsc_clken),
      .line_buf1_Ix_rsc_q(line_buf1_Ix_rsc_q),
      .line_buf1_Ix_rsc_we(line_buf1_Ix_rsc_we),
      .line_buf1_Ix_rsc_d(line_buf1_Ix_rsc_d),
      .line_buf1_Ix_rsc_adr(line_buf1_Ix_rsc_adr),
      .line_buf0_Ix_rsc_clken(line_buf0_Ix_rsc_clken),
      .line_buf0_Ix_rsc_q(line_buf0_Ix_rsc_q),
      .line_buf0_Ix_rsc_we(line_buf0_Ix_rsc_we),
      .line_buf0_Ix_rsc_d(line_buf0_Ix_rsc_d),
      .line_buf0_Ix_rsc_adr(line_buf0_Ix_rsc_adr),
      .line_buf5_Iy_rsc_clken(line_buf5_Iy_rsc_clken),
      .line_buf5_Iy_rsc_q(line_buf5_Iy_rsc_q),
      .line_buf5_Iy_rsc_we(line_buf5_Iy_rsc_we),
      .line_buf5_Iy_rsc_d(line_buf5_Iy_rsc_d),
      .line_buf5_Iy_rsc_adr(line_buf5_Iy_rsc_adr),
      .line_buf4_Iy_rsc_clken(line_buf4_Iy_rsc_clken),
      .line_buf4_Iy_rsc_q(line_buf4_Iy_rsc_q),
      .line_buf4_Iy_rsc_we(line_buf4_Iy_rsc_we),
      .line_buf4_Iy_rsc_d(line_buf4_Iy_rsc_d),
      .line_buf4_Iy_rsc_adr(line_buf4_Iy_rsc_adr),
      .line_buf3_Iy_rsc_clken(line_buf3_Iy_rsc_clken),
      .line_buf3_Iy_rsc_q(line_buf3_Iy_rsc_q),
      .line_buf3_Iy_rsc_we(line_buf3_Iy_rsc_we),
      .line_buf3_Iy_rsc_d(line_buf3_Iy_rsc_d),
      .line_buf3_Iy_rsc_adr(line_buf3_Iy_rsc_adr),
      .line_buf2_Iy_rsc_clken(line_buf2_Iy_rsc_clken),
      .line_buf2_Iy_rsc_q(line_buf2_Iy_rsc_q),
      .line_buf2_Iy_rsc_we(line_buf2_Iy_rsc_we),
      .line_buf2_Iy_rsc_d(line_buf2_Iy_rsc_d),
      .line_buf2_Iy_rsc_adr(line_buf2_Iy_rsc_adr),
      .line_buf1_Iy_rsc_clken(line_buf1_Iy_rsc_clken),
      .line_buf1_Iy_rsc_q(line_buf1_Iy_rsc_q),
      .line_buf1_Iy_rsc_we(line_buf1_Iy_rsc_we),
      .line_buf1_Iy_rsc_d(line_buf1_Iy_rsc_d),
      .line_buf1_Iy_rsc_adr(line_buf1_Iy_rsc_adr),
      .line_buf0_Iy_rsc_clken(line_buf0_Iy_rsc_clken),
      .line_buf0_Iy_rsc_q(line_buf0_Iy_rsc_q),
      .line_buf0_Iy_rsc_we(line_buf0_Iy_rsc_we),
      .line_buf0_Iy_rsc_d(line_buf0_Iy_rsc_d),
      .line_buf0_Iy_rsc_adr(line_buf0_Iy_rsc_adr),
      .line_buf5_Iz_rsc_clken(line_buf5_Iz_rsc_clken),
      .line_buf5_Iz_rsc_q(line_buf5_Iz_rsc_q),
      .line_buf5_Iz_rsc_we(line_buf5_Iz_rsc_we),
      .line_buf5_Iz_rsc_d(line_buf5_Iz_rsc_d),
      .line_buf5_Iz_rsc_adr(line_buf5_Iz_rsc_adr),
      .line_buf4_Iz_rsc_clken(line_buf4_Iz_rsc_clken),
      .line_buf4_Iz_rsc_q(line_buf4_Iz_rsc_q),
      .line_buf4_Iz_rsc_we(line_buf4_Iz_rsc_we),
      .line_buf4_Iz_rsc_d(line_buf4_Iz_rsc_d),
      .line_buf4_Iz_rsc_adr(line_buf4_Iz_rsc_adr),
      .line_buf3_Iz_rsc_clken(line_buf3_Iz_rsc_clken),
      .line_buf3_Iz_rsc_q(line_buf3_Iz_rsc_q),
      .line_buf3_Iz_rsc_we(line_buf3_Iz_rsc_we),
      .line_buf3_Iz_rsc_d(line_buf3_Iz_rsc_d),
      .line_buf3_Iz_rsc_adr(line_buf3_Iz_rsc_adr),
      .line_buf2_Iz_rsc_clken(line_buf2_Iz_rsc_clken),
      .line_buf2_Iz_rsc_q(line_buf2_Iz_rsc_q),
      .line_buf2_Iz_rsc_we(line_buf2_Iz_rsc_we),
      .line_buf2_Iz_rsc_d(line_buf2_Iz_rsc_d),
      .line_buf2_Iz_rsc_adr(line_buf2_Iz_rsc_adr),
      .line_buf1_Iz_rsc_clken(line_buf1_Iz_rsc_clken),
      .line_buf1_Iz_rsc_q(line_buf1_Iz_rsc_q),
      .line_buf1_Iz_rsc_we(line_buf1_Iz_rsc_we),
      .line_buf1_Iz_rsc_d(line_buf1_Iz_rsc_d),
      .line_buf1_Iz_rsc_adr(line_buf1_Iz_rsc_adr),
      .line_buf0_Iz_rsc_clken(line_buf0_Iz_rsc_clken),
      .line_buf0_Iz_rsc_q(line_buf0_Iz_rsc_q),
      .line_buf0_Iz_rsc_we(line_buf0_Iz_rsc_we),
      .line_buf0_Iz_rsc_d(line_buf0_Iz_rsc_d),
      .line_buf0_Iz_rsc_adr(line_buf0_Iz_rsc_adr)
    );
  assign y_filtered_rsc_dat = {y_filtered_rsc_dat_z , y_filtered_rsc_dat_y , y_filtered_rsc_dat_x};
endmodule




//------> ../OpticalFlow_gradient_z_calc.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Sun Jun 16 20:58:56 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_z_calc_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module OpticalFlow_gradient_z_calc_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for OpticalFlow_gradient_z_calc_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : OpticalFlow_gradient_z_calc_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_z_calc_run_staller
// ------------------------------------------------------------------


module OpticalFlow_gradient_z_calc_run_staller (
  run_wen, input_frames_delayed_rsci_wen_comp, gradient_z_rsci_wen_comp
);
  output run_wen;
  input input_frames_delayed_rsci_wen_comp;
  input gradient_z_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = input_frames_delayed_rsci_wen_comp & gradient_z_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_z_calc_run_gradient_z_rsci_gradient_z_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_gradient_z_calc_run_gradient_z_rsci_gradient_z_wait_dp (
  clk, rst, arst_n, gradient_z_rsci_oswt, gradient_z_rsci_wen_comp, gradient_z_rsci_biwt,
      gradient_z_rsci_bdwt, gradient_z_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input gradient_z_rsci_oswt;
  output gradient_z_rsci_wen_comp;
  input gradient_z_rsci_biwt;
  input gradient_z_rsci_bdwt;
  output gradient_z_rsci_bcwt;
  reg gradient_z_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign gradient_z_rsci_wen_comp = (~ gradient_z_rsci_oswt) | gradient_z_rsci_biwt
      | gradient_z_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      gradient_z_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      gradient_z_rsci_bcwt <= 1'b0;
    end
    else begin
      gradient_z_rsci_bcwt <= ~((~(gradient_z_rsci_bcwt | gradient_z_rsci_biwt))
          | gradient_z_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_z_calc_run_gradient_z_rsci_gradient_z_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_z_calc_run_gradient_z_rsci_gradient_z_wait_ctrl (
  run_wen, gradient_z_rsci_oswt, gradient_z_rsci_biwt, gradient_z_rsci_bdwt, gradient_z_rsci_bcwt,
      gradient_z_rsci_irdy, gradient_z_rsci_ivld_run_sct
);
  input run_wen;
  input gradient_z_rsci_oswt;
  output gradient_z_rsci_biwt;
  output gradient_z_rsci_bdwt;
  input gradient_z_rsci_bcwt;
  input gradient_z_rsci_irdy;
  output gradient_z_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire gradient_z_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign gradient_z_rsci_bdwt = gradient_z_rsci_oswt & run_wen;
  assign gradient_z_rsci_biwt = gradient_z_rsci_ogwt & gradient_z_rsci_irdy;
  assign gradient_z_rsci_ogwt = gradient_z_rsci_oswt & (~ gradient_z_rsci_bcwt);
  assign gradient_z_rsci_ivld_run_sct = gradient_z_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_z_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_z_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_ctrl
    (
  run_wen, input_frames_delayed_rsci_iswt0, input_frames_delayed_rsci_irdy_run_sct
);
  input run_wen;
  input input_frames_delayed_rsci_iswt0;
  output input_frames_delayed_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign input_frames_delayed_rsci_irdy_run_sct = input_frames_delayed_rsci_iswt0
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_z_calc_run_gradient_z_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_z_calc_run_gradient_z_rsci (
  clk, rst, arst_n, gradient_z_rsc_dat, gradient_z_rsc_vld, gradient_z_rsc_rdy, run_wen,
      gradient_z_rsci_oswt, gradient_z_rsci_wen_comp, gradient_z_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [31:0] gradient_z_rsc_dat;
  output gradient_z_rsc_vld;
  input gradient_z_rsc_rdy;
  input run_wen;
  input gradient_z_rsci_oswt;
  output gradient_z_rsci_wen_comp;
  input [31:0] gradient_z_rsci_idat;


  // Interconnect Declarations
  wire gradient_z_rsci_biwt;
  wire gradient_z_rsci_bdwt;
  wire gradient_z_rsci_bcwt;
  wire gradient_z_rsci_irdy;
  wire gradient_z_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd32)) gradient_z_rsci (
      .irdy(gradient_z_rsci_irdy),
      .ivld(gradient_z_rsci_ivld_run_sct),
      .idat(gradient_z_rsci_idat),
      .rdy(gradient_z_rsc_rdy),
      .vld(gradient_z_rsc_vld),
      .dat(gradient_z_rsc_dat)
    );
  OpticalFlow_gradient_z_calc_run_gradient_z_rsci_gradient_z_wait_ctrl OpticalFlow_gradient_z_calc_run_gradient_z_rsci_gradient_z_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .gradient_z_rsci_oswt(gradient_z_rsci_oswt),
      .gradient_z_rsci_biwt(gradient_z_rsci_biwt),
      .gradient_z_rsci_bdwt(gradient_z_rsci_bdwt),
      .gradient_z_rsci_bcwt(gradient_z_rsci_bcwt),
      .gradient_z_rsci_irdy(gradient_z_rsci_irdy),
      .gradient_z_rsci_ivld_run_sct(gradient_z_rsci_ivld_run_sct)
    );
  OpticalFlow_gradient_z_calc_run_gradient_z_rsci_gradient_z_wait_dp OpticalFlow_gradient_z_calc_run_gradient_z_rsci_gradient_z_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .gradient_z_rsci_oswt(gradient_z_rsci_oswt),
      .gradient_z_rsci_wen_comp(gradient_z_rsci_wen_comp),
      .gradient_z_rsci_biwt(gradient_z_rsci_biwt),
      .gradient_z_rsci_bdwt(gradient_z_rsci_bdwt),
      .gradient_z_rsci_bcwt(gradient_z_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_z_calc_run_input_frames_delayed_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_z_calc_run_input_frames_delayed_rsci (
  input_frames_delayed_rsc_dat, input_frames_delayed_rsc_vld, input_frames_delayed_rsc_rdy,
      run_wen, input_frames_delayed_rsci_oswt, input_frames_delayed_rsci_wen_comp,
      input_frames_delayed_rsci_idat_mxwt
);
  input [31:0] input_frames_delayed_rsc_dat;
  input input_frames_delayed_rsc_vld;
  output input_frames_delayed_rsc_rdy;
  input run_wen;
  input input_frames_delayed_rsci_oswt;
  output input_frames_delayed_rsci_wen_comp;
  output [31:0] input_frames_delayed_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_frames_delayed_rsci_irdy_run_sct;
  wire input_frames_delayed_rsci_ivld;
  wire [31:0] input_frames_delayed_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd1),
  .width(32'sd32)) input_frames_delayed_rsci (
      .rdy(input_frames_delayed_rsc_rdy),
      .vld(input_frames_delayed_rsc_vld),
      .dat(input_frames_delayed_rsc_dat),
      .irdy(input_frames_delayed_rsci_irdy_run_sct),
      .ivld(input_frames_delayed_rsci_ivld),
      .idat(input_frames_delayed_rsci_idat)
    );
  OpticalFlow_gradient_z_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_ctrl
      OpticalFlow_gradient_z_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .input_frames_delayed_rsci_iswt0(input_frames_delayed_rsci_oswt),
      .input_frames_delayed_rsci_irdy_run_sct(input_frames_delayed_rsci_irdy_run_sct)
    );
  assign input_frames_delayed_rsci_idat_mxwt = input_frames_delayed_rsci_idat;
  assign input_frames_delayed_rsci_wen_comp = (~ input_frames_delayed_rsci_oswt)
      | input_frames_delayed_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_z_calc_run
// ------------------------------------------------------------------


module OpticalFlow_gradient_z_calc_run (
  clk, rst, arst_n, input_frames_delayed_rsc_dat, input_frames_delayed_rsc_vld, input_frames_delayed_rsc_rdy,
      gradient_z_rsc_dat, gradient_z_rsc_vld, gradient_z_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] input_frames_delayed_rsc_dat;
  input input_frames_delayed_rsc_vld;
  output input_frames_delayed_rsc_rdy;
  output [31:0] gradient_z_rsc_dat;
  output gradient_z_rsc_vld;
  input gradient_z_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire input_frames_delayed_rsci_wen_comp;
  wire [31:0] input_frames_delayed_rsci_idat_mxwt;
  wire gradient_z_rsci_wen_comp;
  reg [27:0] gradient_z_rsci_idat_27_0;
  wire [1:0] fsm_output;
  reg main_stage_0_3;
  reg reg_gradient_z_rsci_iswt0_cse;
  reg reg_input_frames_delayed_rsci_iswt0_cse;
  reg main_stage_0_2;
  reg [36:0] Gradient_z_calc_COLUMN_mul_2_itm_1;
  reg [34:0] Gradient_z_calc_COLUMN_mul_3_itm_1;
  wire signed [35:0] nl_Gradient_z_calc_COLUMN_mul_3_itm_1;
  reg [33:0] Gradient_z_calc_COLUMN_mul_itm_1;
  reg [37:0] Gradient_z_calc_COLUMN_acc_6_itm_1;
  wire [38:0] nl_Gradient_z_calc_COLUMN_acc_6_itm_1;
  reg [37:0] Gradient_z_calc_COLUMN_mul_1_itm_1;
  wire signed [38:0] nl_Gradient_z_calc_COLUMN_mul_1_itm_1;
  reg [37:0] Gradient_z_calc_COLUMN_mul_1_itm_2;

  wire[37:0] Gradient_z_calc_COLUMN_acc_nl;
  wire[38:0] nl_Gradient_z_calc_COLUMN_acc_nl;
  wire[34:0] Gradient_z_calc_COLUMN_acc_5_nl;
  wire[35:0] nl_Gradient_z_calc_COLUMN_acc_5_nl;
  wire[24:0] Gradient_z_calc_COLUMN_acc_7_nl;
  wire[25:0] nl_Gradient_z_calc_COLUMN_acc_7_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_OpticalFlow_gradient_z_calc_run_gradient_z_rsci_inst_gradient_z_rsci_idat;
  assign nl_OpticalFlow_gradient_z_calc_run_gradient_z_rsci_inst_gradient_z_rsci_idat
      = {{4{gradient_z_rsci_idat_27_0[27]}}, gradient_z_rsci_idat_27_0};
  OpticalFlow_gradient_z_calc_run_input_frames_delayed_rsci OpticalFlow_gradient_z_calc_run_input_frames_delayed_rsci_inst
      (
      .input_frames_delayed_rsc_dat(input_frames_delayed_rsc_dat),
      .input_frames_delayed_rsc_vld(input_frames_delayed_rsc_vld),
      .input_frames_delayed_rsc_rdy(input_frames_delayed_rsc_rdy),
      .run_wen(run_wen),
      .input_frames_delayed_rsci_oswt(reg_input_frames_delayed_rsci_iswt0_cse),
      .input_frames_delayed_rsci_wen_comp(input_frames_delayed_rsci_wen_comp),
      .input_frames_delayed_rsci_idat_mxwt(input_frames_delayed_rsci_idat_mxwt)
    );
  OpticalFlow_gradient_z_calc_run_gradient_z_rsci OpticalFlow_gradient_z_calc_run_gradient_z_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .gradient_z_rsc_dat(gradient_z_rsc_dat),
      .gradient_z_rsc_vld(gradient_z_rsc_vld),
      .gradient_z_rsc_rdy(gradient_z_rsc_rdy),
      .run_wen(run_wen),
      .gradient_z_rsci_oswt(reg_gradient_z_rsci_iswt0_cse),
      .gradient_z_rsci_wen_comp(gradient_z_rsci_wen_comp),
      .gradient_z_rsci_idat(nl_OpticalFlow_gradient_z_calc_run_gradient_z_rsci_inst_gradient_z_rsci_idat[31:0])
    );
  OpticalFlow_gradient_z_calc_run_staller OpticalFlow_gradient_z_calc_run_staller_inst
      (
      .run_wen(run_wen),
      .input_frames_delayed_rsci_wen_comp(input_frames_delayed_rsci_wen_comp),
      .gradient_z_rsci_wen_comp(gradient_z_rsci_wen_comp)
    );
  OpticalFlow_gradient_z_calc_run_run_fsm OpticalFlow_gradient_z_calc_run_run_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      gradient_z_rsci_idat_27_0 <= 28'b0000000000000000000000000000;
    end
    else if ( rst ) begin
      gradient_z_rsci_idat_27_0 <= 28'b0000000000000000000000000000;
    end
    else if ( run_wen & main_stage_0_3 ) begin
      gradient_z_rsci_idat_27_0 <= readslicef_38_28_10(Gradient_z_calc_COLUMN_acc_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_gradient_z_rsci_iswt0_cse <= 1'b0;
      reg_input_frames_delayed_rsci_iswt0_cse <= 1'b0;
      Gradient_z_calc_COLUMN_acc_6_itm_1 <= 38'b00000000000000000000000000000000000000;
      Gradient_z_calc_COLUMN_mul_1_itm_2 <= 38'b00000000000000000000000000000000000000;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      Gradient_z_calc_COLUMN_mul_2_itm_1 <= 37'b0000000000000000000000000000000000000;
      Gradient_z_calc_COLUMN_mul_3_itm_1 <= 35'b00000000000000000000000000000000000;
      Gradient_z_calc_COLUMN_mul_itm_1 <= 34'b0000000000000000000000000000000000;
      Gradient_z_calc_COLUMN_mul_1_itm_1 <= 38'b00000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      reg_gradient_z_rsci_iswt0_cse <= 1'b0;
      reg_input_frames_delayed_rsci_iswt0_cse <= 1'b0;
      Gradient_z_calc_COLUMN_acc_6_itm_1 <= 38'b00000000000000000000000000000000000000;
      Gradient_z_calc_COLUMN_mul_1_itm_2 <= 38'b00000000000000000000000000000000000000;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      Gradient_z_calc_COLUMN_mul_2_itm_1 <= 37'b0000000000000000000000000000000000000;
      Gradient_z_calc_COLUMN_mul_3_itm_1 <= 35'b00000000000000000000000000000000000;
      Gradient_z_calc_COLUMN_mul_itm_1 <= 34'b0000000000000000000000000000000000;
      Gradient_z_calc_COLUMN_mul_1_itm_1 <= 38'b00000000000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_gradient_z_rsci_iswt0_cse <= main_stage_0_3;
      reg_input_frames_delayed_rsci_iswt0_cse <= 1'b1;
      Gradient_z_calc_COLUMN_acc_6_itm_1 <= nl_Gradient_z_calc_COLUMN_acc_6_itm_1[37:0];
      Gradient_z_calc_COLUMN_mul_1_itm_2 <= Gradient_z_calc_COLUMN_mul_1_itm_1;
      main_stage_0_2 <= fsm_output[1];
      main_stage_0_3 <= main_stage_0_2;
      Gradient_z_calc_COLUMN_mul_2_itm_1 <= (input_frames_delayed_rsci_idat_mxwt[23:16])
          * 29'b10101010101011001101100111101;
      Gradient_z_calc_COLUMN_mul_3_itm_1 <= nl_Gradient_z_calc_COLUMN_mul_3_itm_1[34:0];
      Gradient_z_calc_COLUMN_mul_itm_1 <= (input_frames_delayed_rsci_idat_mxwt[7:0])
          * 26'b10101010100110010011000011;
      Gradient_z_calc_COLUMN_mul_1_itm_1 <= nl_Gradient_z_calc_COLUMN_mul_1_itm_1[37:0];
    end
  end
  assign nl_Gradient_z_calc_COLUMN_acc_nl = Gradient_z_calc_COLUMN_acc_6_itm_1 +
      Gradient_z_calc_COLUMN_mul_1_itm_2;
  assign Gradient_z_calc_COLUMN_acc_nl = nl_Gradient_z_calc_COLUMN_acc_nl[37:0];
  assign nl_Gradient_z_calc_COLUMN_acc_7_nl = (Gradient_z_calc_COLUMN_mul_itm_1[33:9])
      + 25'b0000000000000000000000001;
  assign Gradient_z_calc_COLUMN_acc_7_nl = nl_Gradient_z_calc_COLUMN_acc_7_nl[24:0];
  assign nl_Gradient_z_calc_COLUMN_acc_5_nl = Gradient_z_calc_COLUMN_mul_3_itm_1
      + conv_u2s_34_35({Gradient_z_calc_COLUMN_acc_7_nl , (Gradient_z_calc_COLUMN_mul_itm_1[8:0])});
  assign Gradient_z_calc_COLUMN_acc_5_nl = nl_Gradient_z_calc_COLUMN_acc_5_nl[34:0];
  assign nl_Gradient_z_calc_COLUMN_acc_6_itm_1  = conv_u2s_37_38(Gradient_z_calc_COLUMN_mul_2_itm_1)
      + conv_s2s_35_38(Gradient_z_calc_COLUMN_acc_5_nl);
  assign nl_Gradient_z_calc_COLUMN_mul_3_itm_1  = $signed(conv_u2s_8_9(input_frames_delayed_rsci_idat_mxwt[31:24]))
      * $signed(27'b101010101011001101100111101);
  assign nl_Gradient_z_calc_COLUMN_mul_1_itm_1  = $signed(conv_u2s_8_9(input_frames_delayed_rsci_idat_mxwt[15:8]))
      * $signed(30'b101010101010100110010011000011);

  function automatic [27:0] readslicef_38_28_10;
    input [37:0] vector;
    reg [37:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_38_28_10 = tmp[27:0];
  end
  endfunction


  function automatic [37:0] conv_s2s_35_38 ;
    input [34:0]  vector ;
  begin
    conv_s2s_35_38 = {{3{vector[34]}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [34:0] conv_u2s_34_35 ;
    input [33:0]  vector ;
  begin
    conv_u2s_34_35 =  {1'b0, vector};
  end
  endfunction


  function automatic [37:0] conv_u2s_37_38 ;
    input [36:0]  vector ;
  begin
    conv_u2s_37_38 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_z_calc
// ------------------------------------------------------------------


module OpticalFlow_gradient_z_calc (
  clk, rst, arst_n, input_frames_delayed_rsc_dat, input_frames_delayed_rsc_vld, input_frames_delayed_rsc_rdy,
      gradient_z_rsc_dat, gradient_z_rsc_vld, gradient_z_rsc_rdy, widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] input_frames_delayed_rsc_dat;
  input input_frames_delayed_rsc_vld;
  output input_frames_delayed_rsc_rdy;
  output [31:0] gradient_z_rsc_dat;
  output gradient_z_rsc_vld;
  input gradient_z_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;



  // Interconnect Declarations for Component Instantiations 
  OpticalFlow_gradient_z_calc_run OpticalFlow_gradient_z_calc_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .input_frames_delayed_rsc_dat(input_frames_delayed_rsc_dat),
      .input_frames_delayed_rsc_vld(input_frames_delayed_rsc_vld),
      .input_frames_delayed_rsc_rdy(input_frames_delayed_rsc_rdy),
      .gradient_z_rsc_dat(gradient_z_rsc_dat),
      .gradient_z_rsc_vld(gradient_z_rsc_vld),
      .gradient_z_rsc_rdy(gradient_z_rsc_rdy)
    );
endmodule




//------> ../OpticalFlow_gradient_y_calc.v2/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Sun Jun 16 20:56:47 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_10_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_10_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_9_9_64_512_1_512_64_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_9_9_64_512_1_512_64_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_8_9_16_512_1_512_16_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_8_9_16_512_1_512_16_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [15:0] q;
  output we;
  output [15:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [15:0] d_d;
  output [15:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_7_9_16_512_1_512_16_1_gen
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_7_9_16_512_1_512_16_1_gen
    (
  clken, q, we, d, adr, adr_d, clken_d, d_d, q_d, we_d, rw_rw_ram_ir_internal_RMASK_B_d,
      rw_rw_ram_ir_internal_WMASK_B_d
);
  output clken;
  input [15:0] q;
  output we;
  output [15:0] d;
  output [8:0] adr;
  input [8:0] adr_d;
  input clken_d;
  input [15:0] d_d;
  output [15:0] q_d;
  input we_d;
  input rw_rw_ram_ir_internal_RMASK_B_d;
  input rw_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign we = (rw_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_staller
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_staller (
  run_wen, input_frames_rsci_wen_comp, gradient_y_rsci_wen_comp, frame3_rsci_wen_comp,
      input_frames_delayed_rsci_wen_comp
);
  output run_wen;
  input input_frames_rsci_wen_comp;
  input gradient_y_rsci_wen_comp;
  input frame3_rsci_wen_comp;
  input input_frames_delayed_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = input_frames_rsci_wen_comp & gradient_y_rsci_wen_comp & frame3_rsci_wen_comp
      & input_frames_delayed_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_dp
    (
  clk, rst, arst_n, input_frames_delayed_rsci_oswt, input_frames_delayed_rsci_wen_comp,
      input_frames_delayed_rsci_biwt, input_frames_delayed_rsci_bdwt, input_frames_delayed_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input input_frames_delayed_rsci_oswt;
  output input_frames_delayed_rsci_wen_comp;
  input input_frames_delayed_rsci_biwt;
  input input_frames_delayed_rsci_bdwt;
  output input_frames_delayed_rsci_bcwt;
  reg input_frames_delayed_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign input_frames_delayed_rsci_wen_comp = (~ input_frames_delayed_rsci_oswt)
      | input_frames_delayed_rsci_biwt | input_frames_delayed_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_frames_delayed_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      input_frames_delayed_rsci_bcwt <= 1'b0;
    end
    else begin
      input_frames_delayed_rsci_bcwt <= ~((~(input_frames_delayed_rsci_bcwt | input_frames_delayed_rsci_biwt))
          | input_frames_delayed_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_ctrl
    (
  run_wen, input_frames_delayed_rsci_oswt, input_frames_delayed_rsci_biwt, input_frames_delayed_rsci_bdwt,
      input_frames_delayed_rsci_bcwt, input_frames_delayed_rsci_irdy, input_frames_delayed_rsci_ivld_run_sct
);
  input run_wen;
  input input_frames_delayed_rsci_oswt;
  output input_frames_delayed_rsci_biwt;
  output input_frames_delayed_rsci_bdwt;
  input input_frames_delayed_rsci_bcwt;
  input input_frames_delayed_rsci_irdy;
  output input_frames_delayed_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire input_frames_delayed_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_frames_delayed_rsci_bdwt = input_frames_delayed_rsci_oswt & run_wen;
  assign input_frames_delayed_rsci_biwt = input_frames_delayed_rsci_ogwt & input_frames_delayed_rsci_irdy;
  assign input_frames_delayed_rsci_ogwt = input_frames_delayed_rsci_oswt & (~ input_frames_delayed_rsci_bcwt);
  assign input_frames_delayed_rsci_ivld_run_sct = input_frames_delayed_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_frame3_rsci_frame3_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_frame3_rsci_frame3_wait_dp (
  clk, rst, arst_n, frame3_rsci_oswt, frame3_rsci_wen_comp, frame3_rsci_biwt, frame3_rsci_bdwt,
      frame3_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input frame3_rsci_oswt;
  output frame3_rsci_wen_comp;
  input frame3_rsci_biwt;
  input frame3_rsci_bdwt;
  output frame3_rsci_bcwt;
  reg frame3_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign frame3_rsci_wen_comp = (~ frame3_rsci_oswt) | frame3_rsci_biwt | frame3_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      frame3_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      frame3_rsci_bcwt <= 1'b0;
    end
    else begin
      frame3_rsci_bcwt <= ~((~(frame3_rsci_bcwt | frame3_rsci_biwt)) | frame3_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_frame3_rsci_frame3_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_frame3_rsci_frame3_wait_ctrl (
  run_wen, frame3_rsci_oswt, frame3_rsci_biwt, frame3_rsci_bdwt, frame3_rsci_bcwt,
      frame3_rsci_irdy, frame3_rsci_ivld_run_sct
);
  input run_wen;
  input frame3_rsci_oswt;
  output frame3_rsci_biwt;
  output frame3_rsci_bdwt;
  input frame3_rsci_bcwt;
  input frame3_rsci_irdy;
  output frame3_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire frame3_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign frame3_rsci_bdwt = frame3_rsci_oswt & run_wen;
  assign frame3_rsci_biwt = frame3_rsci_ogwt & frame3_rsci_irdy;
  assign frame3_rsci_ogwt = frame3_rsci_oswt & (~ frame3_rsci_bcwt);
  assign frame3_rsci_ivld_run_sct = frame3_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_gradient_y_rsci_gradient_y_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_gradient_y_rsci_gradient_y_wait_dp (
  clk, rst, arst_n, gradient_y_rsci_oswt, gradient_y_rsci_wen_comp, gradient_y_rsci_biwt,
      gradient_y_rsci_bdwt, gradient_y_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input gradient_y_rsci_oswt;
  output gradient_y_rsci_wen_comp;
  input gradient_y_rsci_biwt;
  input gradient_y_rsci_bdwt;
  output gradient_y_rsci_bcwt;
  reg gradient_y_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign gradient_y_rsci_wen_comp = (~ gradient_y_rsci_oswt) | gradient_y_rsci_biwt
      | gradient_y_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      gradient_y_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      gradient_y_rsci_bcwt <= 1'b0;
    end
    else begin
      gradient_y_rsci_bcwt <= ~((~(gradient_y_rsci_bcwt | gradient_y_rsci_biwt))
          | gradient_y_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_gradient_y_rsci_gradient_y_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_gradient_y_rsci_gradient_y_wait_ctrl (
  run_wen, gradient_y_rsci_oswt, gradient_y_rsci_biwt, gradient_y_rsci_bdwt, gradient_y_rsci_bcwt,
      gradient_y_rsci_irdy, gradient_y_rsci_ivld_run_sct
);
  input run_wen;
  input gradient_y_rsci_oswt;
  output gradient_y_rsci_biwt;
  output gradient_y_rsci_bdwt;
  input gradient_y_rsci_bcwt;
  input gradient_y_rsci_irdy;
  output gradient_y_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire gradient_y_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign gradient_y_rsci_bdwt = gradient_y_rsci_oswt & run_wen;
  assign gradient_y_rsci_biwt = gradient_y_rsci_ogwt & gradient_y_rsci_irdy;
  assign gradient_y_rsci_ogwt = gradient_y_rsci_oswt & (~ gradient_y_rsci_bcwt);
  assign gradient_y_rsci_ivld_run_sct = gradient_y_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_input_frames_rsci_input_frames_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_input_frames_rsci_input_frames_wait_ctrl (
  run_wen, input_frames_rsci_iswt0, input_frames_rsci_irdy_run_sct
);
  input run_wen;
  input input_frames_rsci_iswt0;
  output input_frames_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign input_frames_rsci_irdy_run_sct = input_frames_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci (
  clk, rst, arst_n, input_frames_delayed_rsc_dat, input_frames_delayed_rsc_vld, input_frames_delayed_rsc_rdy,
      run_wen, input_frames_delayed_rsci_oswt, input_frames_delayed_rsci_wen_comp,
      input_frames_delayed_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [31:0] input_frames_delayed_rsc_dat;
  output input_frames_delayed_rsc_vld;
  input input_frames_delayed_rsc_rdy;
  input run_wen;
  input input_frames_delayed_rsci_oswt;
  output input_frames_delayed_rsci_wen_comp;
  input [31:0] input_frames_delayed_rsci_idat;


  // Interconnect Declarations
  wire input_frames_delayed_rsci_biwt;
  wire input_frames_delayed_rsci_bdwt;
  wire input_frames_delayed_rsci_bcwt;
  wire input_frames_delayed_rsci_irdy;
  wire input_frames_delayed_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd32)) input_frames_delayed_rsci (
      .irdy(input_frames_delayed_rsci_irdy),
      .ivld(input_frames_delayed_rsci_ivld_run_sct),
      .idat(input_frames_delayed_rsci_idat),
      .rdy(input_frames_delayed_rsc_rdy),
      .vld(input_frames_delayed_rsc_vld),
      .dat(input_frames_delayed_rsc_dat)
    );
  OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_ctrl
      OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .input_frames_delayed_rsci_oswt(input_frames_delayed_rsci_oswt),
      .input_frames_delayed_rsci_biwt(input_frames_delayed_rsci_biwt),
      .input_frames_delayed_rsci_bdwt(input_frames_delayed_rsci_bdwt),
      .input_frames_delayed_rsci_bcwt(input_frames_delayed_rsci_bcwt),
      .input_frames_delayed_rsci_irdy(input_frames_delayed_rsci_irdy),
      .input_frames_delayed_rsci_ivld_run_sct(input_frames_delayed_rsci_ivld_run_sct)
    );
  OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_dp
      OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci_input_frames_delayed_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .input_frames_delayed_rsci_oswt(input_frames_delayed_rsci_oswt),
      .input_frames_delayed_rsci_wen_comp(input_frames_delayed_rsci_wen_comp),
      .input_frames_delayed_rsci_biwt(input_frames_delayed_rsci_biwt),
      .input_frames_delayed_rsci_bdwt(input_frames_delayed_rsci_bdwt),
      .input_frames_delayed_rsci_bcwt(input_frames_delayed_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_frame3_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_frame3_rsci (
  clk, rst, arst_n, frame3_rsc_dat, frame3_rsc_vld, frame3_rsc_rdy, run_wen, frame3_rsci_oswt,
      frame3_rsci_wen_comp, frame3_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [7:0] frame3_rsc_dat;
  output frame3_rsc_vld;
  input frame3_rsc_rdy;
  input run_wen;
  input frame3_rsci_oswt;
  output frame3_rsci_wen_comp;
  input [7:0] frame3_rsci_idat;


  // Interconnect Declarations
  wire frame3_rsci_biwt;
  wire frame3_rsci_bdwt;
  wire frame3_rsci_bcwt;
  wire frame3_rsci_irdy;
  wire frame3_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd8)) frame3_rsci (
      .irdy(frame3_rsci_irdy),
      .ivld(frame3_rsci_ivld_run_sct),
      .idat(frame3_rsci_idat),
      .rdy(frame3_rsc_rdy),
      .vld(frame3_rsc_vld),
      .dat(frame3_rsc_dat)
    );
  OpticalFlow_gradient_y_calc_run_frame3_rsci_frame3_wait_ctrl OpticalFlow_gradient_y_calc_run_frame3_rsci_frame3_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .frame3_rsci_oswt(frame3_rsci_oswt),
      .frame3_rsci_biwt(frame3_rsci_biwt),
      .frame3_rsci_bdwt(frame3_rsci_bdwt),
      .frame3_rsci_bcwt(frame3_rsci_bcwt),
      .frame3_rsci_irdy(frame3_rsci_irdy),
      .frame3_rsci_ivld_run_sct(frame3_rsci_ivld_run_sct)
    );
  OpticalFlow_gradient_y_calc_run_frame3_rsci_frame3_wait_dp OpticalFlow_gradient_y_calc_run_frame3_rsci_frame3_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .frame3_rsci_oswt(frame3_rsci_oswt),
      .frame3_rsci_wen_comp(frame3_rsci_wen_comp),
      .frame3_rsci_biwt(frame3_rsci_biwt),
      .frame3_rsci_bdwt(frame3_rsci_bdwt),
      .frame3_rsci_bcwt(frame3_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_gradient_y_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_gradient_y_rsci (
  clk, rst, arst_n, gradient_y_rsc_dat, gradient_y_rsc_vld, gradient_y_rsc_rdy, run_wen,
      gradient_y_rsci_oswt, gradient_y_rsci_wen_comp, gradient_y_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [31:0] gradient_y_rsc_dat;
  output gradient_y_rsc_vld;
  input gradient_y_rsc_rdy;
  input run_wen;
  input gradient_y_rsci_oswt;
  output gradient_y_rsci_wen_comp;
  input [31:0] gradient_y_rsci_idat;


  // Interconnect Declarations
  wire gradient_y_rsci_biwt;
  wire gradient_y_rsci_bdwt;
  wire gradient_y_rsci_bcwt;
  wire gradient_y_rsci_irdy;
  wire gradient_y_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd32)) gradient_y_rsci (
      .irdy(gradient_y_rsci_irdy),
      .ivld(gradient_y_rsci_ivld_run_sct),
      .idat(gradient_y_rsci_idat),
      .rdy(gradient_y_rsc_rdy),
      .vld(gradient_y_rsc_vld),
      .dat(gradient_y_rsc_dat)
    );
  OpticalFlow_gradient_y_calc_run_gradient_y_rsci_gradient_y_wait_ctrl OpticalFlow_gradient_y_calc_run_gradient_y_rsci_gradient_y_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .gradient_y_rsci_oswt(gradient_y_rsci_oswt),
      .gradient_y_rsci_biwt(gradient_y_rsci_biwt),
      .gradient_y_rsci_bdwt(gradient_y_rsci_bdwt),
      .gradient_y_rsci_bcwt(gradient_y_rsci_bcwt),
      .gradient_y_rsci_irdy(gradient_y_rsci_irdy),
      .gradient_y_rsci_ivld_run_sct(gradient_y_rsci_ivld_run_sct)
    );
  OpticalFlow_gradient_y_calc_run_gradient_y_rsci_gradient_y_wait_dp OpticalFlow_gradient_y_calc_run_gradient_y_rsci_gradient_y_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .gradient_y_rsci_oswt(gradient_y_rsci_oswt),
      .gradient_y_rsci_wen_comp(gradient_y_rsci_wen_comp),
      .gradient_y_rsci_biwt(gradient_y_rsci_biwt),
      .gradient_y_rsci_bdwt(gradient_y_rsci_bdwt),
      .gradient_y_rsci_bcwt(gradient_y_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run_input_frames_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run_input_frames_rsci (
  input_frames_rsc_dat, input_frames_rsc_vld, input_frames_rsc_rdy, run_wen, input_frames_rsci_oswt,
      input_frames_rsci_wen_comp, input_frames_rsci_idat_mxwt
);
  input [31:0] input_frames_rsc_dat;
  input input_frames_rsc_vld;
  output input_frames_rsc_rdy;
  input run_wen;
  input input_frames_rsci_oswt;
  output input_frames_rsci_wen_comp;
  output [31:0] input_frames_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_frames_rsci_irdy_run_sct;
  wire input_frames_rsci_ivld;
  wire [31:0] input_frames_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd1),
  .width(32'sd32)) input_frames_rsci (
      .rdy(input_frames_rsc_rdy),
      .vld(input_frames_rsc_vld),
      .dat(input_frames_rsc_dat),
      .irdy(input_frames_rsci_irdy_run_sct),
      .ivld(input_frames_rsci_ivld),
      .idat(input_frames_rsci_idat)
    );
  OpticalFlow_gradient_y_calc_run_input_frames_rsci_input_frames_wait_ctrl OpticalFlow_gradient_y_calc_run_input_frames_rsci_input_frames_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .input_frames_rsci_iswt0(input_frames_rsci_oswt),
      .input_frames_rsci_irdy_run_sct(input_frames_rsci_irdy_run_sct)
    );
  assign input_frames_rsci_idat_mxwt = input_frames_rsci_idat;
  assign input_frames_rsci_wen_comp = (~ input_frames_rsci_oswt) | input_frames_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc_run
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc_run (
  clk, rst, arst_n, input_frames_rsc_dat, input_frames_rsc_vld, input_frames_rsc_rdy,
      gradient_y_rsc_dat, gradient_y_rsc_vld, gradient_y_rsc_rdy, frame3_rsc_dat,
      frame3_rsc_vld, frame3_rsc_rdy, input_frames_delayed_rsc_dat, input_frames_delayed_rsc_vld,
      input_frames_delayed_rsc_rdy, widthIn, heightIn, line_buf3_rsci_clken_d, line_buf3_rsci_d_d,
      line_buf3_rsci_q_d, line_buf2_rsci_d_d, line_buf2_rsci_q_d, line_buf1_rsci_d_d,
      line_buf1_rsci_q_d, line_buf0_rsci_d_d, line_buf0_rsci_q_d, line_buf3_rsci_adr_d_pff,
      line_buf3_rsci_we_d_pff, line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] input_frames_rsc_dat;
  input input_frames_rsc_vld;
  output input_frames_rsc_rdy;
  output [31:0] gradient_y_rsc_dat;
  output gradient_y_rsc_vld;
  input gradient_y_rsc_rdy;
  output [7:0] frame3_rsc_dat;
  output frame3_rsc_vld;
  input frame3_rsc_rdy;
  output [31:0] input_frames_delayed_rsc_dat;
  output input_frames_delayed_rsc_vld;
  input input_frames_delayed_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  output line_buf3_rsci_clken_d;
  output [15:0] line_buf3_rsci_d_d;
  input [15:0] line_buf3_rsci_q_d;
  output [15:0] line_buf2_rsci_d_d;
  input [15:0] line_buf2_rsci_q_d;
  output [63:0] line_buf1_rsci_d_d;
  input [63:0] line_buf1_rsci_q_d;
  output [63:0] line_buf0_rsci_d_d;
  input [63:0] line_buf0_rsci_q_d;
  output [8:0] line_buf3_rsci_adr_d_pff;
  output line_buf3_rsci_we_d_pff;
  output line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire input_frames_rsci_wen_comp;
  wire [31:0] input_frames_rsci_idat_mxwt;
  wire gradient_y_rsci_wen_comp;
  wire frame3_rsci_wen_comp;
  reg [7:0] frame3_rsci_idat;
  wire input_frames_delayed_rsci_wen_comp;
  reg [31:0] input_frames_delayed_rsci_idat;
  reg [27:0] gradient_y_rsci_idat_27_0;
  wire [9:0] operator_9_false_acc_tmp;
  wire [10:0] nl_operator_9_false_acc_tmp;
  wire or_dcpl_7;
  wire or_dcpl_8;
  wire and_dcpl_25;
  reg Gradient_y_calc_COLUMN_Gradient_y_calc_COLUMN_if_4_Gradient_y_calc_COLUMN_if_4_nor_svs_1;
  reg operator_9_false_slc_operator_9_false_acc_7_svs_2;
  wire exitL_exit_Gradient_y_calc_ROW_sva_mx0;
  reg operator_9_false_1_slc_operator_9_false_1_acc_8_itm_1;
  reg Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_1;
  reg main_stage_0_4;
  reg [9:0] Gradient_y_calc_COLUMN_x_lpi_1_dfm_1_9_0;
  reg main_stage_0_2;
  reg main_stage_0_3;
  reg operator_9_false_slc_operator_9_false_acc_7_svs_st_1;
  reg main_stage_0_5;
  reg Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_2;
  reg operator_9_false_1_slc_operator_9_false_1_acc_8_itm_2;
  reg Gradient_y_calc_COLUMN_if_slc_Gradient_y_calc_COLUMN_acc_9_svs_1;
  reg Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0;
  wire [8:0] Gradient_y_calc_ROW_y_lpi_1_dfm_1;
  wire exit_Gradient_y_calc_ROW_sva_2_mx0w0;
  reg [10:0] Gradient_y_calc_COLUMN_x_sva_2_1;
  wire [11:0] nl_Gradient_y_calc_COLUMN_x_sva_2_1;
  reg reg_input_frames_delayed_rsci_oswt_cse;
  wire Gradient_y_calc_COLUMN_if_3_and_cse;
  reg reg_input_frames_rsci_oswt_cse;
  wire rdbuf2_pix_and_cse;
  reg [31:0] wrbuf0_pix_31_0_lpi_1_dfm_2;
  wire [31:0] rdbuf1_pix_lpi_1_dfm_1_63_32_mx0;
  wire [7:0] rdbuf1_pix_lpi_1_dfm_1_23_16_2;
  reg [7:0] Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1;
  reg [31:0] input_frames_value_lpi_1_dfm_2;
  reg [15:0] rdbuf2_pix_lpi_1_dfm_1;
  reg [63:0] rdbuf0_pix_lpi_1_dfm_1;
  reg [8:0] Gradient_y_calc_ROW_y_lpi_1_dfm_1_1;
  reg [8:0] Gradient_y_calc_ROW_y_lpi_1_dfm_2;
  reg [7:0] Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_dfm_1;
  reg [7:0] Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_1;
  reg [7:0] Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_2;
  reg [31:0] Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_1;
  reg [31:0] Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_2;
  reg [7:0] Gradient_y_calc_COLUMN_mux_9_itm_1;
  reg [36:0] Gradient_y_calc_COLUMN_mul_1_itm_1;
  reg [34:0] Gradient_y_calc_COLUMN_mul_itm_1;
  wire signed [35:0] nl_Gradient_y_calc_COLUMN_mul_itm_1;
  reg [34:0] Gradient_y_calc_COLUMN_mul_itm_2;
  reg [7:0] Gradient_y_calc_COLUMN_mux_6_itm_1;
  reg [7:0] Gradient_y_calc_COLUMN_mux_7_itm_1;
  reg [37:0] Gradient_y_calc_COLUMN_mul_3_itm_1;
  wire signed [38:0] nl_Gradient_y_calc_COLUMN_mul_3_itm_1;
  reg [7:0] rdbuf3_pix_lpi_1_15_8;
  reg [31:0] rdbuf1_pix_lpi_1_63_32;
  reg [7:0] rdbuf3_pix_lpi_1_dfm_1_15_8;
  reg [31:0] rdbuf1_pix_lpi_1_dfm_1_63_32;
  reg [7:0] rdbuf1_pix_lpi_1_dfm_1_23_16_1;
  reg [7:0] rdbuf2_pix_lpi_1_15_8;
  reg [7:0] rdbuf0_pix_lpi_1_55_48;
  reg [24:0] Gradient_y_calc_COLUMN_acc_6_itm_1_33_9;
  wire [25:0] nl_Gradient_y_calc_COLUMN_acc_6_itm_1_33_9;
  reg [8:0] Gradient_y_calc_COLUMN_acc_6_itm_1_8_0;
  wire gradient_y_rsci_idat_27_0_mx0c1;
  wire [10:0] Gradient_y_calc_COLUMN_x_lpi_1_dfm_2;
  wire [11:0] operator_11_false_acc_psp_sva_1;
  wire [12:0] nl_operator_11_false_acc_psp_sva_1;
  wire [33:0] Gradient_y_calc_COLUMN_mul_4_sdt_1;
  wire [7:0] Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_mx0;
  wire [15:0] rdbuf2_pix_lpi_1_dfm_3;
  wire [31:0] wrbuf0_pix_31_0_lpi_1_dfm_4;
  wire [63:0] rdbuf0_pix_lpi_1_dfm_3;
  wire operator_9_false_acc_itm_9_1;

  wire[37:0] Gradient_y_calc_COLUMN_acc_nl;
  wire[38:0] nl_Gradient_y_calc_COLUMN_acc_nl;
  wire[37:0] Gradient_y_calc_COLUMN_acc_8_nl;
  wire[38:0] nl_Gradient_y_calc_COLUMN_acc_8_nl;
  wire[34:0] Gradient_y_calc_COLUMN_acc_7_nl;
  wire[35:0] nl_Gradient_y_calc_COLUMN_acc_7_nl;
  wire Gradient_y_calc_COLUMN_if_3_not_1_nl;
  wire[9:0] Gradient_y_calc_COLUMN_aelse_acc_nl;
  wire[10:0] nl_Gradient_y_calc_COLUMN_aelse_acc_nl;
  wire[8:0] operator_9_false_1_acc_nl;
  wire[9:0] nl_operator_9_false_1_acc_nl;
  wire[7:0] operator_9_false_acc_nl;
  wire[8:0] nl_operator_9_false_acc_nl;
  wire[10:0] Gradient_y_calc_COLUMN_if_4_mux_nl;
  wire Gradient_y_calc_ROW_Gradient_y_calc_ROW_Gradient_y_calc_ROW_Gradient_y_calc_ROW_not_nl;
  wire[8:0] Gradient_y_calc_COLUMN_if_4_mux_1_nl;
  wire[8:0] Gradient_y_calc_ROW_acc_nl;
  wire[9:0] nl_Gradient_y_calc_ROW_acc_nl;
  wire Gradient_y_calc_ROW_not_15_nl;
  wire[9:0] operator_9_false_acc_nl_1;
  wire[10:0] nl_operator_9_false_acc_nl_1;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_OpticalFlow_gradient_y_calc_run_gradient_y_rsci_inst_gradient_y_rsci_idat;
  assign nl_OpticalFlow_gradient_y_calc_run_gradient_y_rsci_inst_gradient_y_rsci_idat
      = {{4{gradient_y_rsci_idat_27_0[27]}}, gradient_y_rsci_idat_27_0};
  OpticalFlow_gradient_y_calc_run_input_frames_rsci OpticalFlow_gradient_y_calc_run_input_frames_rsci_inst
      (
      .input_frames_rsc_dat(input_frames_rsc_dat),
      .input_frames_rsc_vld(input_frames_rsc_vld),
      .input_frames_rsc_rdy(input_frames_rsc_rdy),
      .run_wen(run_wen),
      .input_frames_rsci_oswt(reg_input_frames_rsci_oswt_cse),
      .input_frames_rsci_wen_comp(input_frames_rsci_wen_comp),
      .input_frames_rsci_idat_mxwt(input_frames_rsci_idat_mxwt)
    );
  OpticalFlow_gradient_y_calc_run_gradient_y_rsci OpticalFlow_gradient_y_calc_run_gradient_y_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .gradient_y_rsc_dat(gradient_y_rsc_dat),
      .gradient_y_rsc_vld(gradient_y_rsc_vld),
      .gradient_y_rsc_rdy(gradient_y_rsc_rdy),
      .run_wen(run_wen),
      .gradient_y_rsci_oswt(reg_input_frames_delayed_rsci_oswt_cse),
      .gradient_y_rsci_wen_comp(gradient_y_rsci_wen_comp),
      .gradient_y_rsci_idat(nl_OpticalFlow_gradient_y_calc_run_gradient_y_rsci_inst_gradient_y_rsci_idat[31:0])
    );
  OpticalFlow_gradient_y_calc_run_frame3_rsci OpticalFlow_gradient_y_calc_run_frame3_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .frame3_rsc_dat(frame3_rsc_dat),
      .frame3_rsc_vld(frame3_rsc_vld),
      .frame3_rsc_rdy(frame3_rsc_rdy),
      .run_wen(run_wen),
      .frame3_rsci_oswt(reg_input_frames_delayed_rsci_oswt_cse),
      .frame3_rsci_wen_comp(frame3_rsci_wen_comp),
      .frame3_rsci_idat(frame3_rsci_idat)
    );
  OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci OpticalFlow_gradient_y_calc_run_input_frames_delayed_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .input_frames_delayed_rsc_dat(input_frames_delayed_rsc_dat),
      .input_frames_delayed_rsc_vld(input_frames_delayed_rsc_vld),
      .input_frames_delayed_rsc_rdy(input_frames_delayed_rsc_rdy),
      .run_wen(run_wen),
      .input_frames_delayed_rsci_oswt(reg_input_frames_delayed_rsci_oswt_cse),
      .input_frames_delayed_rsci_wen_comp(input_frames_delayed_rsci_wen_comp),
      .input_frames_delayed_rsci_idat(input_frames_delayed_rsci_idat)
    );
  OpticalFlow_gradient_y_calc_run_staller OpticalFlow_gradient_y_calc_run_staller_inst
      (
      .run_wen(run_wen),
      .input_frames_rsci_wen_comp(input_frames_rsci_wen_comp),
      .gradient_y_rsci_wen_comp(gradient_y_rsci_wen_comp),
      .frame3_rsci_wen_comp(frame3_rsci_wen_comp),
      .input_frames_delayed_rsci_wen_comp(input_frames_delayed_rsci_wen_comp)
    );
  assign line_buf3_rsci_clken_d = run_wen;
  assign Gradient_y_calc_COLUMN_if_3_and_cse = run_wen & (~ or_dcpl_7);
  assign rdbuf0_pix_lpi_1_dfm_3 = MUX_v_64_2_2(line_buf0_rsci_q_d, rdbuf0_pix_lpi_1_dfm_1,
      or_dcpl_8);
  assign rdbuf2_pix_lpi_1_dfm_3 = MUX_v_16_2_2(line_buf2_rsci_q_d, rdbuf2_pix_lpi_1_dfm_1,
      or_dcpl_8);
  assign wrbuf0_pix_31_0_lpi_1_dfm_4 = MUX_v_32_2_2(input_frames_rsci_idat_mxwt,
      input_frames_value_lpi_1_dfm_2, Gradient_y_calc_COLUMN_if_slc_Gradient_y_calc_COLUMN_acc_9_svs_1);
  assign rdbuf2_pix_and_cse = run_wen & main_stage_0_3;
  assign rdbuf1_pix_lpi_1_dfm_1_63_32_mx0 = MUX_v_32_2_2((line_buf1_rsci_q_d[63:32]),
      rdbuf1_pix_lpi_1_dfm_1_63_32, or_dcpl_8);
  assign rdbuf1_pix_lpi_1_dfm_1_23_16_2 = MUX_v_8_2_2((line_buf1_rsci_q_d[23:16]),
      rdbuf1_pix_lpi_1_dfm_1_23_16_1, or_dcpl_8);
  assign exitL_exit_Gradient_y_calc_ROW_sva_mx0 = ~((~(exit_Gradient_y_calc_ROW_sva_2_mx0w0
      & Gradient_y_calc_COLUMN_Gradient_y_calc_COLUMN_if_4_Gradient_y_calc_COLUMN_if_4_nor_svs_1))
      & main_stage_0_2);
  assign Gradient_y_calc_COLUMN_if_4_mux_nl = MUX_v_11_2_2(Gradient_y_calc_COLUMN_x_sva_2_1,
      ({{10{exit_Gradient_y_calc_ROW_sva_2_mx0w0}}, exit_Gradient_y_calc_ROW_sva_2_mx0w0}),
      Gradient_y_calc_COLUMN_Gradient_y_calc_COLUMN_if_4_Gradient_y_calc_COLUMN_if_4_nor_svs_1);
  assign Gradient_y_calc_ROW_Gradient_y_calc_ROW_Gradient_y_calc_ROW_Gradient_y_calc_ROW_not_nl
      = ~ exitL_exit_Gradient_y_calc_ROW_sva_mx0;
  assign Gradient_y_calc_COLUMN_x_lpi_1_dfm_2 = MUX_v_11_2_2(11'b00000000000, Gradient_y_calc_COLUMN_if_4_mux_nl,
      Gradient_y_calc_ROW_Gradient_y_calc_ROW_Gradient_y_calc_ROW_Gradient_y_calc_ROW_not_nl);
  assign exit_Gradient_y_calc_ROW_sva_2_mx0w0 = ~((Gradient_y_calc_ROW_y_lpi_1_dfm_1_1
      != (operator_9_false_acc_tmp[8:0])) | (operator_9_false_acc_tmp[9]));
  assign nl_Gradient_y_calc_ROW_acc_nl = Gradient_y_calc_ROW_y_lpi_1_dfm_1_1 + 9'b000000001;
  assign Gradient_y_calc_ROW_acc_nl = nl_Gradient_y_calc_ROW_acc_nl[8:0];
  assign Gradient_y_calc_COLUMN_if_4_mux_1_nl = MUX_v_9_2_2(Gradient_y_calc_ROW_y_lpi_1_dfm_1_1,
      Gradient_y_calc_ROW_acc_nl, Gradient_y_calc_COLUMN_Gradient_y_calc_COLUMN_if_4_Gradient_y_calc_COLUMN_if_4_nor_svs_1);
  assign Gradient_y_calc_ROW_not_15_nl = ~ exitL_exit_Gradient_y_calc_ROW_sva_mx0;
  assign Gradient_y_calc_ROW_y_lpi_1_dfm_1 = MUX_v_9_2_2(9'b000000000, Gradient_y_calc_COLUMN_if_4_mux_1_nl,
      Gradient_y_calc_ROW_not_15_nl);
  assign nl_operator_9_false_acc_tmp = conv_u2s_9_10(heightIn) + 10'b0000000001;
  assign operator_9_false_acc_tmp = nl_operator_9_false_acc_tmp[9:0];
  assign nl_operator_9_false_acc_nl_1 = ({1'b1 , heightIn}) + conv_u2s_9_10(~ Gradient_y_calc_ROW_y_lpi_1_dfm_1);
  assign operator_9_false_acc_nl_1 = nl_operator_9_false_acc_nl_1[9:0];
  assign operator_9_false_acc_itm_9_1 = readslicef_10_1_9(operator_9_false_acc_nl_1);
  assign nl_operator_11_false_acc_psp_sva_1 = conv_u2s_11_12(widthIn) + 12'b111111111111;
  assign operator_11_false_acc_psp_sva_1 = nl_operator_11_false_acc_psp_sva_1[11:0];
  assign Gradient_y_calc_COLUMN_mul_4_sdt_1 = Gradient_y_calc_COLUMN_mux_6_itm_1
      * 26'b10101010100110010011000011;
  assign Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_mx0 = MUX_v_8_2_2(Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1,
      Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_dfm_1, main_stage_0_3);
  assign or_dcpl_7 = ~((~((~ Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_2)
      & operator_9_false_1_slc_operator_9_false_1_acc_8_itm_2)) & main_stage_0_5);
  assign or_dcpl_8 = (~ main_stage_0_3) | Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0;
  assign and_dcpl_25 = main_stage_0_3 & (~ Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0);
  assign gradient_y_rsci_idat_27_0_mx0c1 = main_stage_0_5 & (~ Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_2)
      & (~ operator_9_false_1_slc_operator_9_false_1_acc_8_itm_2);
  assign line_buf3_rsci_adr_d_pff = Gradient_y_calc_COLUMN_x_lpi_1_dfm_1_9_0[9:1];
  assign line_buf3_rsci_d_d = rdbuf2_pix_lpi_1_dfm_3;
  assign line_buf3_rsci_we_d_pff = main_stage_0_2 & (Gradient_y_calc_COLUMN_x_lpi_1_dfm_1_9_0[0]);
  assign line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff = ~((~ main_stage_0_2)
      | (Gradient_y_calc_COLUMN_x_lpi_1_dfm_1_9_0[0]));
  assign line_buf2_rsci_d_d = {(rdbuf1_pix_lpi_1_dfm_1_63_32_mx0[23:16]) , rdbuf1_pix_lpi_1_dfm_1_23_16_2};
  assign line_buf1_rsci_d_d = rdbuf0_pix_lpi_1_dfm_3;
  assign line_buf0_rsci_d_d = {wrbuf0_pix_31_0_lpi_1_dfm_4 , wrbuf0_pix_31_0_lpi_1_dfm_2};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_input_frames_delayed_rsci_oswt_cse <= 1'b0;
      Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_2 <= 8'b00000000;
      Gradient_y_calc_COLUMN_mul_1_itm_1 <= 37'b0000000000000000000000000000000000000;
      Gradient_y_calc_COLUMN_mul_itm_2 <= 35'b00000000000000000000000000000000000;
      Gradient_y_calc_COLUMN_acc_6_itm_1_33_9 <= 25'b0000000000000000000000000;
      Gradient_y_calc_COLUMN_acc_6_itm_1_8_0 <= 9'b000000000;
      Gradient_y_calc_COLUMN_mul_3_itm_1 <= 38'b00000000000000000000000000000000000000;
      operator_9_false_1_slc_operator_9_false_1_acc_8_itm_2 <= 1'b0;
      Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_2 <= 1'b0;
      Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_1 <= 1'b0;
      rdbuf1_pix_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf1_pix_lpi_1_dfm_1_23_16_1 <= 8'b00000000;
      rdbuf0_pix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf2_pix_lpi_1_dfm_1 <= 16'b0000000000000000;
      Gradient_y_calc_ROW_y_lpi_1_dfm_2 <= 9'b000000000;
      operator_9_false_slc_operator_9_false_acc_7_svs_2 <= 1'b0;
      Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0 <= 1'b0;
      Gradient_y_calc_COLUMN_x_lpi_1_dfm_1_9_0 <= 10'b0000000000;
      Gradient_y_calc_COLUMN_Gradient_y_calc_COLUMN_if_4_Gradient_y_calc_COLUMN_if_4_nor_svs_1
          <= 1'b0;
      Gradient_y_calc_ROW_y_lpi_1_dfm_1_1 <= 9'b000000000;
      Gradient_y_calc_COLUMN_x_sva_2_1 <= 11'b00000000000;
      Gradient_y_calc_COLUMN_if_slc_Gradient_y_calc_COLUMN_acc_9_svs_1 <= 1'b0;
      reg_input_frames_rsci_oswt_cse <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      Gradient_y_calc_COLUMN_mux_7_itm_1 <= 8'b00000000;
      Gradient_y_calc_COLUMN_mux_6_itm_1 <= 8'b00000000;
      Gradient_y_calc_COLUMN_mux_9_itm_1 <= 8'b00000000;
      operator_9_false_1_slc_operator_9_false_1_acc_8_itm_1 <= 1'b0;
      operator_9_false_slc_operator_9_false_acc_7_svs_st_1 <= 1'b0;
      Gradient_y_calc_COLUMN_mul_itm_1 <= 35'b00000000000000000000000000000000000;
      Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_1 <= 8'b00000000;
      Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_dfm_1 <= 8'b00000000;
      Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1 <= 8'b00000000;
    end
    else if ( rst ) begin
      reg_input_frames_delayed_rsci_oswt_cse <= 1'b0;
      Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
      Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_2 <= 8'b00000000;
      Gradient_y_calc_COLUMN_mul_1_itm_1 <= 37'b0000000000000000000000000000000000000;
      Gradient_y_calc_COLUMN_mul_itm_2 <= 35'b00000000000000000000000000000000000;
      Gradient_y_calc_COLUMN_acc_6_itm_1_33_9 <= 25'b0000000000000000000000000;
      Gradient_y_calc_COLUMN_acc_6_itm_1_8_0 <= 9'b000000000;
      Gradient_y_calc_COLUMN_mul_3_itm_1 <= 38'b00000000000000000000000000000000000000;
      operator_9_false_1_slc_operator_9_false_1_acc_8_itm_2 <= 1'b0;
      Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_2 <= 1'b0;
      Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_1 <= 1'b0;
      rdbuf1_pix_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
      rdbuf1_pix_lpi_1_dfm_1_23_16_1 <= 8'b00000000;
      rdbuf0_pix_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rdbuf2_pix_lpi_1_dfm_1 <= 16'b0000000000000000;
      Gradient_y_calc_ROW_y_lpi_1_dfm_2 <= 9'b000000000;
      operator_9_false_slc_operator_9_false_acc_7_svs_2 <= 1'b0;
      Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0 <= 1'b0;
      Gradient_y_calc_COLUMN_x_lpi_1_dfm_1_9_0 <= 10'b0000000000;
      Gradient_y_calc_COLUMN_Gradient_y_calc_COLUMN_if_4_Gradient_y_calc_COLUMN_if_4_nor_svs_1
          <= 1'b0;
      Gradient_y_calc_ROW_y_lpi_1_dfm_1_1 <= 9'b000000000;
      Gradient_y_calc_COLUMN_x_sva_2_1 <= 11'b00000000000;
      Gradient_y_calc_COLUMN_if_slc_Gradient_y_calc_COLUMN_acc_9_svs_1 <= 1'b0;
      reg_input_frames_rsci_oswt_cse <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      Gradient_y_calc_COLUMN_mux_7_itm_1 <= 8'b00000000;
      Gradient_y_calc_COLUMN_mux_6_itm_1 <= 8'b00000000;
      Gradient_y_calc_COLUMN_mux_9_itm_1 <= 8'b00000000;
      operator_9_false_1_slc_operator_9_false_1_acc_8_itm_1 <= 1'b0;
      operator_9_false_slc_operator_9_false_acc_7_svs_st_1 <= 1'b0;
      Gradient_y_calc_COLUMN_mul_itm_1 <= 35'b00000000000000000000000000000000000;
      Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_1 <= 8'b00000000;
      Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_dfm_1 <= 8'b00000000;
      Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1 <= 8'b00000000;
    end
    else if ( run_wen ) begin
      reg_input_frames_delayed_rsci_oswt_cse <= ~ or_dcpl_7;
      Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_2 <= Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_1;
      Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_2 <= Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_1;
      Gradient_y_calc_COLUMN_mul_1_itm_1 <= Gradient_y_calc_COLUMN_mux_9_itm_1 *
          29'b10101010101011001101100111101;
      Gradient_y_calc_COLUMN_mul_itm_2 <= Gradient_y_calc_COLUMN_mul_itm_1;
      Gradient_y_calc_COLUMN_acc_6_itm_1_33_9 <= nl_Gradient_y_calc_COLUMN_acc_6_itm_1_33_9[24:0];
      Gradient_y_calc_COLUMN_acc_6_itm_1_8_0 <= Gradient_y_calc_COLUMN_mul_4_sdt_1[8:0];
      Gradient_y_calc_COLUMN_mul_3_itm_1 <= nl_Gradient_y_calc_COLUMN_mul_3_itm_1[37:0];
      operator_9_false_1_slc_operator_9_false_1_acc_8_itm_2 <= operator_9_false_1_slc_operator_9_false_1_acc_8_itm_1;
      Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_2 <= Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_1;
      Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_1 <= (readslicef_10_1_9(Gradient_y_calc_COLUMN_aelse_acc_nl))
          & (~ operator_9_false_slc_operator_9_false_acc_7_svs_2);
      rdbuf1_pix_lpi_1_dfm_1_63_32 <= rdbuf1_pix_lpi_1_dfm_1_63_32_mx0;
      rdbuf1_pix_lpi_1_dfm_1_23_16_1 <= rdbuf1_pix_lpi_1_dfm_1_23_16_2;
      rdbuf0_pix_lpi_1_dfm_1 <= rdbuf0_pix_lpi_1_dfm_3;
      rdbuf2_pix_lpi_1_dfm_1 <= rdbuf2_pix_lpi_1_dfm_3;
      Gradient_y_calc_ROW_y_lpi_1_dfm_2 <= Gradient_y_calc_ROW_y_lpi_1_dfm_1_1;
      operator_9_false_slc_operator_9_false_acc_7_svs_2 <= operator_9_false_slc_operator_9_false_acc_7_svs_st_1;
      Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0 <= Gradient_y_calc_COLUMN_x_lpi_1_dfm_1_9_0[0];
      Gradient_y_calc_COLUMN_x_lpi_1_dfm_1_9_0 <= Gradient_y_calc_COLUMN_x_lpi_1_dfm_2[9:0];
      Gradient_y_calc_COLUMN_Gradient_y_calc_COLUMN_if_4_Gradient_y_calc_COLUMN_if_4_nor_svs_1
          <= ~((Gradient_y_calc_COLUMN_x_lpi_1_dfm_2 != (operator_11_false_acc_psp_sva_1[10:0]))
          | (operator_11_false_acc_psp_sva_1[11]));
      Gradient_y_calc_ROW_y_lpi_1_dfm_1_1 <= Gradient_y_calc_ROW_y_lpi_1_dfm_1;
      Gradient_y_calc_COLUMN_x_sva_2_1 <= nl_Gradient_y_calc_COLUMN_x_sva_2_1[10:0];
      Gradient_y_calc_COLUMN_if_slc_Gradient_y_calc_COLUMN_acc_9_svs_1 <= operator_9_false_acc_itm_9_1;
      reg_input_frames_rsci_oswt_cse <= ~ operator_9_false_acc_itm_9_1;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      Gradient_y_calc_COLUMN_mux_7_itm_1 <= MUX_v_8_2_2((line_buf2_rsci_q_d[7:0]),
          rdbuf2_pix_lpi_1_15_8, Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_y_calc_COLUMN_mux_6_itm_1 <= MUX_v_8_2_2((line_buf3_rsci_q_d[7:0]),
          rdbuf3_pix_lpi_1_15_8, Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_y_calc_COLUMN_mux_9_itm_1 <= MUX_v_8_2_2((line_buf0_rsci_q_d[23:16]),
          rdbuf0_pix_lpi_1_55_48, Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0);
      operator_9_false_1_slc_operator_9_false_1_acc_8_itm_1 <= readslicef_9_1_8(operator_9_false_1_acc_nl);
      operator_9_false_slc_operator_9_false_acc_7_svs_st_1 <= readslicef_8_1_7(operator_9_false_acc_nl);
      Gradient_y_calc_COLUMN_mul_itm_1 <= nl_Gradient_y_calc_COLUMN_mul_itm_1[34:0];
      Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_1 <= MUX_v_32_2_2((line_buf1_rsci_q_d[31:0]),
          rdbuf1_pix_lpi_1_63_32, Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_1 <= MUX_v_8_2_2((line_buf1_rsci_q_d[23:16]),
          (rdbuf1_pix_lpi_1_63_32[23:16]), Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0);
      Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_dfm_1 <= MUX_v_8_2_2((input_frames_rsci_idat_mxwt[23:16]),
          Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_mx0, Gradient_y_calc_COLUMN_if_slc_Gradient_y_calc_COLUMN_acc_9_svs_1);
      Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1 <= Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_frames_delayed_rsci_idat <= 32'b00000000000000000000000000000000;
      frame3_rsci_idat <= 8'b00000000;
    end
    else if ( rst ) begin
      input_frames_delayed_rsci_idat <= 32'b00000000000000000000000000000000;
      frame3_rsci_idat <= 8'b00000000;
    end
    else if ( Gradient_y_calc_COLUMN_if_3_and_cse ) begin
      input_frames_delayed_rsci_idat <= Gradient_y_calc_COLUMN_qr_4_lpi_1_dfm_2;
      frame3_rsci_idat <= Gradient_y_calc_COLUMN_qr_2_lpi_1_dfm_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      gradient_y_rsci_idat_27_0 <= 28'b0000000000000000000000000000;
    end
    else if ( rst ) begin
      gradient_y_rsci_idat_27_0 <= 28'b0000000000000000000000000000;
    end
    else if ( run_wen & ((main_stage_0_5 & Gradient_y_calc_COLUMN_if_3_Gradient_y_calc_COLUMN_if_3_and_itm_2)
        | gradient_y_rsci_idat_27_0_mx0c1) ) begin
      gradient_y_rsci_idat_27_0 <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (readslicef_38_28_10(Gradient_y_calc_COLUMN_acc_nl)), Gradient_y_calc_COLUMN_if_3_not_1_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_frames_value_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      input_frames_value_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & (~((~ main_stage_0_2) | Gradient_y_calc_COLUMN_if_slc_Gradient_y_calc_COLUMN_acc_9_svs_1))
        ) begin
      input_frames_value_lpi_1_dfm_2 <= input_frames_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      wrbuf0_pix_31_0_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      wrbuf0_pix_31_0_lpi_1_dfm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & (~ (Gradient_y_calc_COLUMN_x_lpi_1_dfm_1_9_0[0])) ) begin
      wrbuf0_pix_31_0_lpi_1_dfm_2 <= wrbuf0_pix_31_0_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rdbuf2_pix_lpi_1_15_8 <= 8'b00000000;
      rdbuf3_pix_lpi_1_15_8 <= 8'b00000000;
      rdbuf0_pix_lpi_1_55_48 <= 8'b00000000;
      rdbuf1_pix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      rdbuf2_pix_lpi_1_15_8 <= 8'b00000000;
      rdbuf3_pix_lpi_1_15_8 <= 8'b00000000;
      rdbuf0_pix_lpi_1_55_48 <= 8'b00000000;
      rdbuf1_pix_lpi_1_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( rdbuf2_pix_and_cse ) begin
      rdbuf2_pix_lpi_1_15_8 <= MUX_v_8_2_2((line_buf2_rsci_q_d[15:8]), (rdbuf2_pix_lpi_1_dfm_1[15:8]),
          Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf3_pix_lpi_1_15_8 <= MUX_v_8_2_2(rdbuf3_pix_lpi_1_dfm_1_15_8, (line_buf3_rsci_q_d[15:8]),
          and_dcpl_25);
      rdbuf0_pix_lpi_1_55_48 <= MUX_v_8_2_2((line_buf0_rsci_q_d[55:48]), (rdbuf0_pix_lpi_1_dfm_1[55:48]),
          Gradient_y_calc_COLUMN_x_lpi_1_dfm_2_0);
      rdbuf1_pix_lpi_1_63_32 <= MUX_v_32_2_2(rdbuf1_pix_lpi_1_dfm_1_63_32, (line_buf1_rsci_q_d[63:32]),
          and_dcpl_25);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rdbuf3_pix_lpi_1_dfm_1_15_8 <= 8'b00000000;
    end
    else if ( rst ) begin
      rdbuf3_pix_lpi_1_dfm_1_15_8 <= 8'b00000000;
    end
    else if ( run_wen & (~ or_dcpl_8) ) begin
      rdbuf3_pix_lpi_1_dfm_1_15_8 <= line_buf3_rsci_q_d[15:8];
    end
  end
  assign nl_Gradient_y_calc_COLUMN_acc_6_itm_1_33_9  = (Gradient_y_calc_COLUMN_mul_4_sdt_1[33:9])
      + 25'b0000000000000000000000001;
  assign nl_Gradient_y_calc_COLUMN_mul_3_itm_1  = $signed(conv_u2s_8_9(Gradient_y_calc_COLUMN_mux_7_itm_1))
      * $signed(30'b101010101010100110010011000011);
  assign nl_Gradient_y_calc_COLUMN_aelse_acc_nl = ({1'b1 , Gradient_y_calc_ROW_y_lpi_1_dfm_2})
      + conv_u2u_9_10(~ heightIn) + 10'b0000000001;
  assign Gradient_y_calc_COLUMN_aelse_acc_nl = nl_Gradient_y_calc_COLUMN_aelse_acc_nl[9:0];
  assign nl_Gradient_y_calc_COLUMN_x_sva_2_1  = Gradient_y_calc_COLUMN_x_lpi_1_dfm_2
      + 11'b00000000001;
  assign nl_operator_9_false_1_acc_nl = conv_u2u_8_9(Gradient_y_calc_ROW_y_lpi_1_dfm_2[8:1])
      + 9'b111111111;
  assign operator_9_false_1_acc_nl = nl_operator_9_false_1_acc_nl[8:0];
  assign nl_operator_9_false_acc_nl = conv_u2u_7_8(Gradient_y_calc_ROW_y_lpi_1_dfm_1[8:2])
      + 8'b11111111;
  assign operator_9_false_acc_nl = nl_operator_9_false_acc_nl[7:0];
  assign nl_Gradient_y_calc_COLUMN_mul_itm_1  = $signed(conv_u2s_8_9(Gradient_y_calc_COLUMN_if_ac_fixed_cctor_lpi_1_dfm_1))
      * $signed(27'b101010101011001101100111101);
  assign nl_Gradient_y_calc_COLUMN_acc_7_nl = Gradient_y_calc_COLUMN_mul_itm_2 +
      conv_u2s_34_35({Gradient_y_calc_COLUMN_acc_6_itm_1_33_9 , Gradient_y_calc_COLUMN_acc_6_itm_1_8_0});
  assign Gradient_y_calc_COLUMN_acc_7_nl = nl_Gradient_y_calc_COLUMN_acc_7_nl[34:0];
  assign nl_Gradient_y_calc_COLUMN_acc_8_nl = conv_u2s_37_38(Gradient_y_calc_COLUMN_mul_1_itm_1)
      + conv_s2s_35_38(Gradient_y_calc_COLUMN_acc_7_nl);
  assign Gradient_y_calc_COLUMN_acc_8_nl = nl_Gradient_y_calc_COLUMN_acc_8_nl[37:0];
  assign nl_Gradient_y_calc_COLUMN_acc_nl = Gradient_y_calc_COLUMN_acc_8_nl + Gradient_y_calc_COLUMN_mul_3_itm_1;
  assign Gradient_y_calc_COLUMN_acc_nl = nl_Gradient_y_calc_COLUMN_acc_nl[37:0];
  assign Gradient_y_calc_COLUMN_if_3_not_1_nl = ~ gradient_y_rsci_idat_27_0_mx0c1;

  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [27:0] MUX_v_28_2_2;
    input [27:0] input_0;
    input [27:0] input_1;
    input  sel;
    reg [27:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_28_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [27:0] readslicef_38_28_10;
    input [37:0] vector;
    reg [37:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_38_28_10 = tmp[27:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [37:0] conv_s2s_35_38 ;
    input [34:0]  vector ;
  begin
    conv_s2s_35_38 = {{3{vector[34]}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [34:0] conv_u2s_34_35 ;
    input [33:0]  vector ;
  begin
    conv_u2s_34_35 =  {1'b0, vector};
  end
  endfunction


  function automatic [37:0] conv_u2s_37_38 ;
    input [36:0]  vector ;
  begin
    conv_u2s_37_38 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_y_calc
// ------------------------------------------------------------------


module OpticalFlow_gradient_y_calc (
  clk, rst, arst_n, input_frames_rsc_dat, input_frames_rsc_vld, input_frames_rsc_rdy,
      gradient_y_rsc_dat, gradient_y_rsc_vld, gradient_y_rsc_rdy, frame3_rsc_dat,
      frame3_rsc_vld, frame3_rsc_rdy, input_frames_delayed_rsc_dat, input_frames_delayed_rsc_vld,
      input_frames_delayed_rsc_rdy, widthIn, heightIn, line_buf3_rsc_clken, line_buf3_rsc_q,
      line_buf3_rsc_we, line_buf3_rsc_d, line_buf3_rsc_adr, line_buf2_rsc_clken,
      line_buf2_rsc_q, line_buf2_rsc_we, line_buf2_rsc_d, line_buf2_rsc_adr, line_buf1_rsc_clken,
      line_buf1_rsc_q, line_buf1_rsc_we, line_buf1_rsc_d, line_buf1_rsc_adr, line_buf0_rsc_clken,
      line_buf0_rsc_q, line_buf0_rsc_we, line_buf0_rsc_d, line_buf0_rsc_adr
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] input_frames_rsc_dat;
  input input_frames_rsc_vld;
  output input_frames_rsc_rdy;
  output [31:0] gradient_y_rsc_dat;
  output gradient_y_rsc_vld;
  input gradient_y_rsc_rdy;
  output [7:0] frame3_rsc_dat;
  output frame3_rsc_vld;
  input frame3_rsc_rdy;
  output [31:0] input_frames_delayed_rsc_dat;
  output input_frames_delayed_rsc_vld;
  input input_frames_delayed_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  output line_buf3_rsc_clken;
  input [15:0] line_buf3_rsc_q;
  output line_buf3_rsc_we;
  output [15:0] line_buf3_rsc_d;
  output [8:0] line_buf3_rsc_adr;
  output line_buf2_rsc_clken;
  input [15:0] line_buf2_rsc_q;
  output line_buf2_rsc_we;
  output [15:0] line_buf2_rsc_d;
  output [8:0] line_buf2_rsc_adr;
  output line_buf1_rsc_clken;
  input [63:0] line_buf1_rsc_q;
  output line_buf1_rsc_we;
  output [63:0] line_buf1_rsc_d;
  output [8:0] line_buf1_rsc_adr;
  output line_buf0_rsc_clken;
  input [63:0] line_buf0_rsc_q;
  output line_buf0_rsc_we;
  output [63:0] line_buf0_rsc_d;
  output [8:0] line_buf0_rsc_adr;


  // Interconnect Declarations
  wire line_buf3_rsci_clken_d;
  wire [15:0] line_buf3_rsci_d_d;
  wire [15:0] line_buf3_rsci_q_d;
  wire [15:0] line_buf2_rsci_d_d;
  wire [15:0] line_buf2_rsci_q_d;
  wire [63:0] line_buf1_rsci_d_d;
  wire [63:0] line_buf1_rsci_q_d;
  wire [63:0] line_buf0_rsci_d_d;
  wire [63:0] line_buf0_rsci_q_d;
  wire [8:0] line_buf3_rsci_adr_d_iff;
  wire line_buf3_rsci_we_d_iff;
  wire line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff;


  // Interconnect Declarations for Component Instantiations 
  OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_7_9_16_512_1_512_16_1_gen
      line_buf3_rsci (
      .clken(line_buf3_rsc_clken),
      .q(line_buf3_rsc_q),
      .we(line_buf3_rsc_we),
      .d(line_buf3_rsc_d),
      .adr(line_buf3_rsc_adr),
      .adr_d(line_buf3_rsci_adr_d_iff),
      .clken_d(line_buf3_rsci_clken_d),
      .d_d(line_buf3_rsci_d_d),
      .q_d(line_buf3_rsci_q_d),
      .we_d(line_buf3_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf3_rsci_we_d_iff)
    );
  OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_8_9_16_512_1_512_16_1_gen
      line_buf2_rsci (
      .clken(line_buf2_rsc_clken),
      .q(line_buf2_rsc_q),
      .we(line_buf2_rsc_we),
      .d(line_buf2_rsc_d),
      .adr(line_buf2_rsc_adr),
      .adr_d(line_buf3_rsci_adr_d_iff),
      .clken_d(line_buf3_rsci_clken_d),
      .d_d(line_buf2_rsci_d_d),
      .q_d(line_buf2_rsci_q_d),
      .we_d(line_buf3_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf3_rsci_we_d_iff)
    );
  OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_9_9_64_512_1_512_64_1_gen
      line_buf1_rsci (
      .clken(line_buf1_rsc_clken),
      .q(line_buf1_rsc_q),
      .we(line_buf1_rsc_we),
      .d(line_buf1_rsc_d),
      .adr(line_buf1_rsc_adr),
      .adr_d(line_buf3_rsci_adr_d_iff),
      .clken_d(line_buf3_rsci_clken_d),
      .d_d(line_buf1_rsci_d_d),
      .q_d(line_buf1_rsci_q_d),
      .we_d(line_buf3_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf3_rsci_we_d_iff)
    );
  OpticalFlow_gradient_y_calc_Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_en_10_9_64_512_1_512_64_1_gen
      line_buf0_rsci (
      .clken(line_buf0_rsc_clken),
      .q(line_buf0_rsc_q),
      .we(line_buf0_rsc_we),
      .d(line_buf0_rsc_d),
      .adr(line_buf0_rsc_adr),
      .adr_d(line_buf3_rsci_adr_d_iff),
      .clken_d(line_buf3_rsci_clken_d),
      .d_d(line_buf0_rsci_d_d),
      .q_d(line_buf0_rsci_q_d),
      .we_d(line_buf3_rsci_we_d_iff),
      .rw_rw_ram_ir_internal_RMASK_B_d(line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff),
      .rw_rw_ram_ir_internal_WMASK_B_d(line_buf3_rsci_we_d_iff)
    );
  OpticalFlow_gradient_y_calc_run OpticalFlow_gradient_y_calc_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .input_frames_rsc_dat(input_frames_rsc_dat),
      .input_frames_rsc_vld(input_frames_rsc_vld),
      .input_frames_rsc_rdy(input_frames_rsc_rdy),
      .gradient_y_rsc_dat(gradient_y_rsc_dat),
      .gradient_y_rsc_vld(gradient_y_rsc_vld),
      .gradient_y_rsc_rdy(gradient_y_rsc_rdy),
      .frame3_rsc_dat(frame3_rsc_dat),
      .frame3_rsc_vld(frame3_rsc_vld),
      .frame3_rsc_rdy(frame3_rsc_rdy),
      .input_frames_delayed_rsc_dat(input_frames_delayed_rsc_dat),
      .input_frames_delayed_rsc_vld(input_frames_delayed_rsc_vld),
      .input_frames_delayed_rsc_rdy(input_frames_delayed_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .line_buf3_rsci_clken_d(line_buf3_rsci_clken_d),
      .line_buf3_rsci_d_d(line_buf3_rsci_d_d),
      .line_buf3_rsci_q_d(line_buf3_rsci_q_d),
      .line_buf2_rsci_d_d(line_buf2_rsci_d_d),
      .line_buf2_rsci_q_d(line_buf2_rsci_q_d),
      .line_buf1_rsci_d_d(line_buf1_rsci_d_d),
      .line_buf1_rsci_q_d(line_buf1_rsci_q_d),
      .line_buf0_rsci_d_d(line_buf0_rsci_d_d),
      .line_buf0_rsci_q_d(line_buf0_rsci_q_d),
      .line_buf3_rsci_adr_d_pff(line_buf3_rsci_adr_d_iff),
      .line_buf3_rsci_we_d_pff(line_buf3_rsci_we_d_iff),
      .line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_pff(line_buf3_rsci_rw_rw_ram_ir_internal_RMASK_B_d_iff)
    );
endmodule




//------> ../OpticalFlow_gradient_x_calc.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Sun Jun 16 20:51:51 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_x_calc_run_staller
// ------------------------------------------------------------------


module OpticalFlow_gradient_x_calc_run_staller (
  run_wen, frame3_b_rsci_wen_comp, gradient_x_rsci_wen_comp
);
  output run_wen;
  input frame3_b_rsci_wen_comp;
  input gradient_x_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = frame3_b_rsci_wen_comp & gradient_x_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_x_calc_run_gradient_x_rsci_gradient_x_wait_dp
// ------------------------------------------------------------------


module OpticalFlow_gradient_x_calc_run_gradient_x_rsci_gradient_x_wait_dp (
  clk, rst, arst_n, gradient_x_rsci_oswt, gradient_x_rsci_wen_comp, gradient_x_rsci_biwt,
      gradient_x_rsci_bdwt, gradient_x_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input gradient_x_rsci_oswt;
  output gradient_x_rsci_wen_comp;
  input gradient_x_rsci_biwt;
  input gradient_x_rsci_bdwt;
  output gradient_x_rsci_bcwt;
  reg gradient_x_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign gradient_x_rsci_wen_comp = (~ gradient_x_rsci_oswt) | gradient_x_rsci_biwt
      | gradient_x_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      gradient_x_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      gradient_x_rsci_bcwt <= 1'b0;
    end
    else begin
      gradient_x_rsci_bcwt <= ~((~(gradient_x_rsci_bcwt | gradient_x_rsci_biwt))
          | gradient_x_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_x_calc_run_gradient_x_rsci_gradient_x_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_x_calc_run_gradient_x_rsci_gradient_x_wait_ctrl (
  run_wen, gradient_x_rsci_oswt, gradient_x_rsci_biwt, gradient_x_rsci_bdwt, gradient_x_rsci_bcwt,
      gradient_x_rsci_irdy, gradient_x_rsci_ivld_run_sct
);
  input run_wen;
  input gradient_x_rsci_oswt;
  output gradient_x_rsci_biwt;
  output gradient_x_rsci_bdwt;
  input gradient_x_rsci_bcwt;
  input gradient_x_rsci_irdy;
  output gradient_x_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire gradient_x_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign gradient_x_rsci_bdwt = gradient_x_rsci_oswt & run_wen;
  assign gradient_x_rsci_biwt = gradient_x_rsci_ogwt & gradient_x_rsci_irdy;
  assign gradient_x_rsci_ogwt = gradient_x_rsci_oswt & (~ gradient_x_rsci_bcwt);
  assign gradient_x_rsci_ivld_run_sct = gradient_x_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_x_calc_run_frame3_b_rsci_frame3_b_wait_ctrl
// ------------------------------------------------------------------


module OpticalFlow_gradient_x_calc_run_frame3_b_rsci_frame3_b_wait_ctrl (
  run_wen, frame3_b_rsci_iswt0, frame3_b_rsci_irdy_run_sct
);
  input run_wen;
  input frame3_b_rsci_iswt0;
  output frame3_b_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign frame3_b_rsci_irdy_run_sct = frame3_b_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_x_calc_run_gradient_x_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_x_calc_run_gradient_x_rsci (
  clk, rst, arst_n, gradient_x_rsc_dat, gradient_x_rsc_vld, gradient_x_rsc_rdy, run_wen,
      gradient_x_rsci_oswt, gradient_x_rsci_wen_comp, gradient_x_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [31:0] gradient_x_rsc_dat;
  output gradient_x_rsc_vld;
  input gradient_x_rsc_rdy;
  input run_wen;
  input gradient_x_rsci_oswt;
  output gradient_x_rsci_wen_comp;
  input [31:0] gradient_x_rsci_idat;


  // Interconnect Declarations
  wire gradient_x_rsci_biwt;
  wire gradient_x_rsci_bdwt;
  wire gradient_x_rsci_bcwt;
  wire gradient_x_rsci_irdy;
  wire gradient_x_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd32)) gradient_x_rsci (
      .irdy(gradient_x_rsci_irdy),
      .ivld(gradient_x_rsci_ivld_run_sct),
      .idat(gradient_x_rsci_idat),
      .rdy(gradient_x_rsc_rdy),
      .vld(gradient_x_rsc_vld),
      .dat(gradient_x_rsc_dat)
    );
  OpticalFlow_gradient_x_calc_run_gradient_x_rsci_gradient_x_wait_ctrl OpticalFlow_gradient_x_calc_run_gradient_x_rsci_gradient_x_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .gradient_x_rsci_oswt(gradient_x_rsci_oswt),
      .gradient_x_rsci_biwt(gradient_x_rsci_biwt),
      .gradient_x_rsci_bdwt(gradient_x_rsci_bdwt),
      .gradient_x_rsci_bcwt(gradient_x_rsci_bcwt),
      .gradient_x_rsci_irdy(gradient_x_rsci_irdy),
      .gradient_x_rsci_ivld_run_sct(gradient_x_rsci_ivld_run_sct)
    );
  OpticalFlow_gradient_x_calc_run_gradient_x_rsci_gradient_x_wait_dp OpticalFlow_gradient_x_calc_run_gradient_x_rsci_gradient_x_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .gradient_x_rsci_oswt(gradient_x_rsci_oswt),
      .gradient_x_rsci_wen_comp(gradient_x_rsci_wen_comp),
      .gradient_x_rsci_biwt(gradient_x_rsci_biwt),
      .gradient_x_rsci_bdwt(gradient_x_rsci_bdwt),
      .gradient_x_rsci_bcwt(gradient_x_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_x_calc_run_frame3_b_rsci
// ------------------------------------------------------------------


module OpticalFlow_gradient_x_calc_run_frame3_b_rsci (
  frame3_b_rsc_dat, frame3_b_rsc_vld, frame3_b_rsc_rdy, run_wen, frame3_b_rsci_oswt,
      frame3_b_rsci_wen_comp, frame3_b_rsci_idat_mxwt
);
  input [7:0] frame3_b_rsc_dat;
  input frame3_b_rsc_vld;
  output frame3_b_rsc_rdy;
  input run_wen;
  input frame3_b_rsci_oswt;
  output frame3_b_rsci_wen_comp;
  output [7:0] frame3_b_rsci_idat_mxwt;


  // Interconnect Declarations
  wire frame3_b_rsci_irdy_run_sct;
  wire frame3_b_rsci_ivld;
  wire [7:0] frame3_b_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd1),
  .width(32'sd8)) frame3_b_rsci (
      .rdy(frame3_b_rsc_rdy),
      .vld(frame3_b_rsc_vld),
      .dat(frame3_b_rsc_dat),
      .irdy(frame3_b_rsci_irdy_run_sct),
      .ivld(frame3_b_rsci_ivld),
      .idat(frame3_b_rsci_idat)
    );
  OpticalFlow_gradient_x_calc_run_frame3_b_rsci_frame3_b_wait_ctrl OpticalFlow_gradient_x_calc_run_frame3_b_rsci_frame3_b_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .frame3_b_rsci_iswt0(frame3_b_rsci_oswt),
      .frame3_b_rsci_irdy_run_sct(frame3_b_rsci_irdy_run_sct)
    );
  assign frame3_b_rsci_idat_mxwt = frame3_b_rsci_idat;
  assign frame3_b_rsci_wen_comp = (~ frame3_b_rsci_oswt) | frame3_b_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_x_calc_run
// ------------------------------------------------------------------


module OpticalFlow_gradient_x_calc_run (
  clk, rst, arst_n, frame3_b_rsc_dat, frame3_b_rsc_vld, frame3_b_rsc_rdy, gradient_x_rsc_dat,
      gradient_x_rsc_vld, gradient_x_rsc_rdy, widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [7:0] frame3_b_rsc_dat;
  input frame3_b_rsc_vld;
  output frame3_b_rsc_rdy;
  output [31:0] gradient_x_rsc_dat;
  output gradient_x_rsc_vld;
  input gradient_x_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;


  // Interconnect Declarations
  wire run_wen;
  wire frame3_b_rsci_wen_comp;
  wire [7:0] frame3_b_rsci_idat_mxwt;
  wire gradient_x_rsci_wen_comp;
  reg [27:0] gradient_x_rsci_idat_27_0;
  wire [9:0] operator_9_false_acc_tmp;
  wire [10:0] nl_operator_9_false_acc_tmp;
  wire Gradient_x_calc_COLUMN_Gradient_x_calc_COLUMN_if_2_nor_tmp;
  wire exit_Gradient_x_calc_ROW_sva_2_mx0;
  reg Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_1;
  reg main_stage_0_2;
  reg main_stage_0_3;
  reg Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_2;
  reg operator_11_false_1_slc_operator_11_false_1_acc_10_itm_2;
  reg Gradient_x_calc_COLUMN_if_2_and_itm_1;
  reg Gradient_x_calc_COLUMN_if_slc_Gradient_x_calc_COLUMN_acc_11_svs_1;
  wire [10:0] Gradient_x_calc_COLUMN_x_lpi_1_dfm_3;
  reg reg_gradient_x_rsci_oswt_cse;
  reg reg_frame3_b_rsci_oswt_cse;
  wire [7:0] pix_buf0_mux_cse;
  reg [7:0] pix_buf2_lpi_1;
  reg exitL_exit_Gradient_x_calc_ROW_sva;
  reg exit_Gradient_x_calc_ROW_sva_2;
  reg [10:0] Gradient_x_calc_COLUMN_x_lpi_1_dfm_2;
  reg exit_Gradient_x_calc_ROW_lpi_1_dfm_2;
  reg [8:0] Gradient_x_calc_ROW_y_sva_1_1;
  wire [9:0] nl_Gradient_x_calc_ROW_y_sva_1_1;
  reg [7:0] pix_buf0_lpi_1_dfm_1;
  reg [7:0] pix_buf2_lpi_1_dfm_1;
  reg [8:0] Gradient_x_calc_ROW_y_lpi_1_dfm_1;
  reg [36:0] Gradient_x_calc_COLUMN_mul_1_itm_1;
  reg [34:0] Gradient_x_calc_COLUMN_mul_itm_1;
  wire signed [35:0] nl_Gradient_x_calc_COLUMN_mul_itm_1;
  reg [7:0] Gradient_x_calc_ROW_Gradient_x_calc_ROW_and_3_itm_1;
  reg [37:0] Gradient_x_calc_COLUMN_mul_3_itm_1;
  wire signed [38:0] nl_Gradient_x_calc_COLUMN_mul_3_itm_1;
  reg operator_11_false_1_slc_operator_11_false_1_acc_10_itm_1;
  reg [24:0] Gradient_x_calc_COLUMN_acc_7_itm_1_33_9;
  wire [25:0] nl_Gradient_x_calc_COLUMN_acc_7_itm_1_33_9;
  reg [8:0] Gradient_x_calc_COLUMN_acc_7_itm_1_8_0;
  wire gradient_x_rsci_idat_27_0_mx0c1;
  wire [8:0] Gradient_x_calc_ROW_y_lpi_1_dfm_1_1;
  wire exit_Gradient_x_calc_ROW_sva_2_mx0w0;
  wire [11:0] operator_11_false_return_11_0_sva_1;
  wire [12:0] nl_operator_11_false_return_11_0_sva_1;
  wire exit_Gradient_x_calc_ROW_lpi_1_dfm_3;
  wire [33:0] Gradient_x_calc_COLUMN_mul_4_sdt_1;
  wire operator_11_false_acc_itm_11_1;

  wire[37:0] Gradient_x_calc_COLUMN_acc_nl;
  wire[38:0] nl_Gradient_x_calc_COLUMN_acc_nl;
  wire[37:0] Gradient_x_calc_COLUMN_acc_9_nl;
  wire[38:0] nl_Gradient_x_calc_COLUMN_acc_9_nl;
  wire[34:0] Gradient_x_calc_COLUMN_acc_8_nl;
  wire[35:0] nl_Gradient_x_calc_COLUMN_acc_8_nl;
  wire Gradient_x_calc_COLUMN_if_1_not_2_nl;
  wire[11:0] Gradient_x_calc_COLUMN_aelse_acc_nl;
  wire[12:0] nl_Gradient_x_calc_COLUMN_aelse_acc_nl;
  wire[9:0] operator_11_false_acc_nl;
  wire[10:0] nl_operator_11_false_acc_nl;
  wire[10:0] Gradient_x_calc_COLUMN_acc_5_nl;
  wire[11:0] nl_Gradient_x_calc_COLUMN_acc_5_nl;
  wire Gradient_x_calc_ROW_not_22_nl;
  wire Gradient_x_calc_ROW_not_21_nl;
  wire Gradient_x_calc_ROW_not_23_nl;
  wire[10:0] operator_11_false_1_acc_nl;
  wire[11:0] nl_operator_11_false_1_acc_nl;
  wire Gradient_x_calc_ROW_not_18_nl;
  wire[8:0] Gradient_x_calc_ROW_y_mux_nl;
  wire Gradient_x_calc_ROW_not_20_nl;
  wire[11:0] operator_11_false_acc_nl_1;
  wire[12:0] nl_operator_11_false_acc_nl_1;
  wire Gradient_x_calc_ROW_Gradient_x_calc_ROW_Gradient_x_calc_ROW_nor_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_OpticalFlow_gradient_x_calc_run_gradient_x_rsci_inst_gradient_x_rsci_idat;
  assign nl_OpticalFlow_gradient_x_calc_run_gradient_x_rsci_inst_gradient_x_rsci_idat
      = {{4{gradient_x_rsci_idat_27_0[27]}}, gradient_x_rsci_idat_27_0};
  OpticalFlow_gradient_x_calc_run_frame3_b_rsci OpticalFlow_gradient_x_calc_run_frame3_b_rsci_inst
      (
      .frame3_b_rsc_dat(frame3_b_rsc_dat),
      .frame3_b_rsc_vld(frame3_b_rsc_vld),
      .frame3_b_rsc_rdy(frame3_b_rsc_rdy),
      .run_wen(run_wen),
      .frame3_b_rsci_oswt(reg_frame3_b_rsci_oswt_cse),
      .frame3_b_rsci_wen_comp(frame3_b_rsci_wen_comp),
      .frame3_b_rsci_idat_mxwt(frame3_b_rsci_idat_mxwt)
    );
  OpticalFlow_gradient_x_calc_run_gradient_x_rsci OpticalFlow_gradient_x_calc_run_gradient_x_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .gradient_x_rsc_dat(gradient_x_rsc_dat),
      .gradient_x_rsc_vld(gradient_x_rsc_vld),
      .gradient_x_rsc_rdy(gradient_x_rsc_rdy),
      .run_wen(run_wen),
      .gradient_x_rsci_oswt(reg_gradient_x_rsci_oswt_cse),
      .gradient_x_rsci_wen_comp(gradient_x_rsci_wen_comp),
      .gradient_x_rsci_idat(nl_OpticalFlow_gradient_x_calc_run_gradient_x_rsci_inst_gradient_x_rsci_idat[31:0])
    );
  OpticalFlow_gradient_x_calc_run_staller OpticalFlow_gradient_x_calc_run_staller_inst
      (
      .run_wen(run_wen),
      .frame3_b_rsci_wen_comp(frame3_b_rsci_wen_comp),
      .gradient_x_rsci_wen_comp(gradient_x_rsci_wen_comp)
    );
  assign pix_buf0_mux_cse = MUX_v_8_2_2(frame3_b_rsci_idat_mxwt, pix_buf0_lpi_1_dfm_1,
      Gradient_x_calc_COLUMN_if_slc_Gradient_x_calc_COLUMN_acc_11_svs_1);
  assign Gradient_x_calc_ROW_y_mux_nl = MUX_v_9_2_2(Gradient_x_calc_ROW_y_lpi_1_dfm_1,
      Gradient_x_calc_ROW_y_sva_1_1, Gradient_x_calc_COLUMN_if_2_and_itm_1);
  assign Gradient_x_calc_ROW_not_20_nl = ~ exitL_exit_Gradient_x_calc_ROW_sva;
  assign Gradient_x_calc_ROW_y_lpi_1_dfm_1_1 = MUX_v_9_2_2(9'b000000000, Gradient_x_calc_ROW_y_mux_nl,
      Gradient_x_calc_ROW_not_20_nl);
  assign nl_operator_11_false_acc_nl_1 = ({1'b1 , widthIn}) + conv_u2s_11_12(~ Gradient_x_calc_COLUMN_x_lpi_1_dfm_3);
  assign operator_11_false_acc_nl_1 = nl_operator_11_false_acc_nl_1[11:0];
  assign operator_11_false_acc_itm_11_1 = readslicef_12_1_11(operator_11_false_acc_nl_1);
  assign Gradient_x_calc_ROW_Gradient_x_calc_ROW_Gradient_x_calc_ROW_nor_nl = ~(exit_Gradient_x_calc_ROW_lpi_1_dfm_2
      | exitL_exit_Gradient_x_calc_ROW_sva);
  assign Gradient_x_calc_COLUMN_x_lpi_1_dfm_3 = MUX_v_11_2_2(11'b00000000000, Gradient_x_calc_COLUMN_x_lpi_1_dfm_2,
      Gradient_x_calc_ROW_Gradient_x_calc_ROW_Gradient_x_calc_ROW_nor_nl);
  assign exit_Gradient_x_calc_ROW_sva_2_mx0w0 = ~((Gradient_x_calc_ROW_y_lpi_1_dfm_1_1
      != (operator_9_false_acc_tmp[8:0])) | (operator_9_false_acc_tmp[9]));
  assign exit_Gradient_x_calc_ROW_sva_2_mx0 = MUX_s_1_2_2(exit_Gradient_x_calc_ROW_sva_2,
      exit_Gradient_x_calc_ROW_sva_2_mx0w0, Gradient_x_calc_COLUMN_Gradient_x_calc_COLUMN_if_2_nor_tmp);
  assign nl_operator_9_false_acc_tmp = conv_u2s_9_10(heightIn) + 10'b1111111111;
  assign operator_9_false_acc_tmp = nl_operator_9_false_acc_tmp[9:0];
  assign Gradient_x_calc_COLUMN_Gradient_x_calc_COLUMN_if_2_nor_tmp = ~((Gradient_x_calc_COLUMN_x_lpi_1_dfm_3
      != (operator_11_false_return_11_0_sva_1[10:0])) | (operator_11_false_return_11_0_sva_1[11]));
  assign nl_operator_11_false_return_11_0_sva_1 = conv_u2s_11_12(widthIn) + 12'b000000000001;
  assign operator_11_false_return_11_0_sva_1 = nl_operator_11_false_return_11_0_sva_1[11:0];
  assign exit_Gradient_x_calc_ROW_lpi_1_dfm_3 = exit_Gradient_x_calc_ROW_sva_2_mx0
      & Gradient_x_calc_COLUMN_Gradient_x_calc_COLUMN_if_2_nor_tmp;
  assign Gradient_x_calc_COLUMN_mul_4_sdt_1 = Gradient_x_calc_ROW_Gradient_x_calc_ROW_and_3_itm_1
      * 26'b10101010100110010011000011;
  assign gradient_x_rsci_idat_27_0_mx0c1 = main_stage_0_3 & (~ operator_11_false_1_slc_operator_11_false_1_acc_10_itm_2)
      & (~ Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_2);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_gradient_x_rsci_oswt_cse <= 1'b0;
      Gradient_x_calc_COLUMN_mul_1_itm_1 <= 37'b0000000000000000000000000000000000000;
      Gradient_x_calc_COLUMN_mul_itm_1 <= 35'b00000000000000000000000000000000000;
      Gradient_x_calc_COLUMN_acc_7_itm_1_33_9 <= 25'b0000000000000000000000000;
      Gradient_x_calc_COLUMN_acc_7_itm_1_8_0 <= 9'b000000000;
      Gradient_x_calc_COLUMN_mul_3_itm_1 <= 38'b00000000000000000000000000000000000000;
      operator_11_false_1_slc_operator_11_false_1_acc_10_itm_2 <= 1'b0;
      Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_2 <= 1'b0;
      Gradient_x_calc_ROW_y_lpi_1_dfm_1 <= 9'b000000000;
      Gradient_x_calc_ROW_y_sva_1_1 <= 9'b000000000;
      Gradient_x_calc_COLUMN_if_2_and_itm_1 <= 1'b0;
      Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_1 <= 1'b0;
      reg_frame3_b_rsci_oswt_cse <= 1'b0;
      exit_Gradient_x_calc_ROW_sva_2 <= 1'b0;
      Gradient_x_calc_COLUMN_x_lpi_1_dfm_2 <= 11'b00000000000;
      exit_Gradient_x_calc_ROW_lpi_1_dfm_2 <= 1'b0;
      exitL_exit_Gradient_x_calc_ROW_sva <= 1'b1;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      pix_buf2_lpi_1_dfm_1 <= 8'b00000000;
      Gradient_x_calc_ROW_Gradient_x_calc_ROW_and_3_itm_1 <= 8'b00000000;
      pix_buf0_lpi_1_dfm_1 <= 8'b00000000;
      Gradient_x_calc_COLUMN_if_slc_Gradient_x_calc_COLUMN_acc_11_svs_1 <= 1'b0;
      operator_11_false_1_slc_operator_11_false_1_acc_10_itm_1 <= 1'b0;
      pix_buf2_lpi_1 <= 8'b00000000;
    end
    else if ( rst ) begin
      reg_gradient_x_rsci_oswt_cse <= 1'b0;
      Gradient_x_calc_COLUMN_mul_1_itm_1 <= 37'b0000000000000000000000000000000000000;
      Gradient_x_calc_COLUMN_mul_itm_1 <= 35'b00000000000000000000000000000000000;
      Gradient_x_calc_COLUMN_acc_7_itm_1_33_9 <= 25'b0000000000000000000000000;
      Gradient_x_calc_COLUMN_acc_7_itm_1_8_0 <= 9'b000000000;
      Gradient_x_calc_COLUMN_mul_3_itm_1 <= 38'b00000000000000000000000000000000000000;
      operator_11_false_1_slc_operator_11_false_1_acc_10_itm_2 <= 1'b0;
      Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_2 <= 1'b0;
      Gradient_x_calc_ROW_y_lpi_1_dfm_1 <= 9'b000000000;
      Gradient_x_calc_ROW_y_sva_1_1 <= 9'b000000000;
      Gradient_x_calc_COLUMN_if_2_and_itm_1 <= 1'b0;
      Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_1 <= 1'b0;
      reg_frame3_b_rsci_oswt_cse <= 1'b0;
      exit_Gradient_x_calc_ROW_sva_2 <= 1'b0;
      Gradient_x_calc_COLUMN_x_lpi_1_dfm_2 <= 11'b00000000000;
      exit_Gradient_x_calc_ROW_lpi_1_dfm_2 <= 1'b0;
      exitL_exit_Gradient_x_calc_ROW_sva <= 1'b1;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      pix_buf2_lpi_1_dfm_1 <= 8'b00000000;
      Gradient_x_calc_ROW_Gradient_x_calc_ROW_and_3_itm_1 <= 8'b00000000;
      pix_buf0_lpi_1_dfm_1 <= 8'b00000000;
      Gradient_x_calc_COLUMN_if_slc_Gradient_x_calc_COLUMN_acc_11_svs_1 <= 1'b0;
      operator_11_false_1_slc_operator_11_false_1_acc_10_itm_1 <= 1'b0;
      pix_buf2_lpi_1 <= 8'b00000000;
    end
    else if ( run_wen ) begin
      reg_gradient_x_rsci_oswt_cse <= (~(operator_11_false_1_slc_operator_11_false_1_acc_10_itm_2
          & (~ Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_2)))
          & main_stage_0_3;
      Gradient_x_calc_COLUMN_mul_1_itm_1 <= pix_buf0_lpi_1_dfm_1 * 29'b10101010101011001101100111101;
      Gradient_x_calc_COLUMN_mul_itm_1 <= nl_Gradient_x_calc_COLUMN_mul_itm_1[34:0];
      Gradient_x_calc_COLUMN_acc_7_itm_1_33_9 <= nl_Gradient_x_calc_COLUMN_acc_7_itm_1_33_9[24:0];
      Gradient_x_calc_COLUMN_acc_7_itm_1_8_0 <= Gradient_x_calc_COLUMN_mul_4_sdt_1[8:0];
      Gradient_x_calc_COLUMN_mul_3_itm_1 <= nl_Gradient_x_calc_COLUMN_mul_3_itm_1[37:0];
      operator_11_false_1_slc_operator_11_false_1_acc_10_itm_2 <= operator_11_false_1_slc_operator_11_false_1_acc_10_itm_1;
      Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_2 <= Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_1;
      Gradient_x_calc_ROW_y_lpi_1_dfm_1 <= Gradient_x_calc_ROW_y_lpi_1_dfm_1_1;
      Gradient_x_calc_ROW_y_sva_1_1 <= nl_Gradient_x_calc_ROW_y_sva_1_1[8:0];
      Gradient_x_calc_COLUMN_if_2_and_itm_1 <= (~ exit_Gradient_x_calc_ROW_sva_2_mx0)
          & Gradient_x_calc_COLUMN_Gradient_x_calc_COLUMN_if_2_nor_tmp;
      Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_1 <= (readslicef_12_1_11(Gradient_x_calc_COLUMN_aelse_acc_nl))
          & (~ (readslicef_10_1_9(operator_11_false_acc_nl)));
      reg_frame3_b_rsci_oswt_cse <= ~ operator_11_false_acc_itm_11_1;
      exit_Gradient_x_calc_ROW_sva_2 <= exit_Gradient_x_calc_ROW_sva_2_mx0;
      Gradient_x_calc_COLUMN_x_lpi_1_dfm_2 <= MUX_v_11_2_2(Gradient_x_calc_COLUMN_acc_5_nl,
          ({{10{exit_Gradient_x_calc_ROW_sva_2_mx0w0}}, exit_Gradient_x_calc_ROW_sva_2_mx0w0}),
          Gradient_x_calc_COLUMN_Gradient_x_calc_COLUMN_if_2_nor_tmp);
      exit_Gradient_x_calc_ROW_lpi_1_dfm_2 <= exit_Gradient_x_calc_ROW_lpi_1_dfm_3;
      exitL_exit_Gradient_x_calc_ROW_sva <= exit_Gradient_x_calc_ROW_lpi_1_dfm_3;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      pix_buf2_lpi_1_dfm_1 <= MUX_v_8_2_2(8'b00000000, pix_buf2_lpi_1, Gradient_x_calc_ROW_not_22_nl);
      Gradient_x_calc_ROW_Gradient_x_calc_ROW_and_3_itm_1 <= MUX_v_8_2_2(8'b00000000,
          pix_buf2_lpi_1_dfm_1, Gradient_x_calc_ROW_not_21_nl);
      pix_buf0_lpi_1_dfm_1 <= MUX_v_8_2_2(8'b00000000, pix_buf0_mux_cse, Gradient_x_calc_ROW_not_23_nl);
      Gradient_x_calc_COLUMN_if_slc_Gradient_x_calc_COLUMN_acc_11_svs_1 <= operator_11_false_acc_itm_11_1;
      operator_11_false_1_slc_operator_11_false_1_acc_10_itm_1 <= readslicef_11_1_10(operator_11_false_1_acc_nl);
      pix_buf2_lpi_1 <= MUX_v_8_2_2(8'b00000000, pix_buf0_lpi_1_dfm_1, Gradient_x_calc_ROW_not_18_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      gradient_x_rsci_idat_27_0 <= 28'b0000000000000000000000000000;
    end
    else if ( rst ) begin
      gradient_x_rsci_idat_27_0 <= 28'b0000000000000000000000000000;
    end
    else if ( run_wen & ((main_stage_0_3 & Gradient_x_calc_COLUMN_if_1_Gradient_x_calc_COLUMN_if_1_and_itm_2)
        | gradient_x_rsci_idat_27_0_mx0c1) ) begin
      gradient_x_rsci_idat_27_0 <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (readslicef_38_28_10(Gradient_x_calc_COLUMN_acc_nl)), Gradient_x_calc_COLUMN_if_1_not_2_nl);
    end
  end
  assign nl_Gradient_x_calc_COLUMN_mul_itm_1  = $signed(conv_u2s_8_9(pix_buf0_mux_cse))
      * $signed(27'b101010101011001101100111101);
  assign nl_Gradient_x_calc_COLUMN_acc_7_itm_1_33_9  = (Gradient_x_calc_COLUMN_mul_4_sdt_1[33:9])
      + 25'b0000000000000000000000001;
  assign nl_Gradient_x_calc_COLUMN_mul_3_itm_1  = $signed(conv_u2s_8_9(pix_buf2_lpi_1_dfm_1))
      * $signed(30'b101010101010100110010011000011);
  assign nl_Gradient_x_calc_ROW_y_sva_1_1  = Gradient_x_calc_ROW_y_lpi_1_dfm_1_1
      + 9'b000000001;
  assign nl_Gradient_x_calc_COLUMN_aelse_acc_nl = ({1'b1 , Gradient_x_calc_COLUMN_x_lpi_1_dfm_3})
      + conv_u2u_11_12(~ widthIn) + 12'b000000000001;
  assign Gradient_x_calc_COLUMN_aelse_acc_nl = nl_Gradient_x_calc_COLUMN_aelse_acc_nl[11:0];
  assign nl_operator_11_false_acc_nl = conv_u2u_9_10(Gradient_x_calc_COLUMN_x_lpi_1_dfm_3[10:2])
      + 10'b1111111111;
  assign operator_11_false_acc_nl = nl_operator_11_false_acc_nl[9:0];
  assign nl_Gradient_x_calc_COLUMN_acc_5_nl = Gradient_x_calc_COLUMN_x_lpi_1_dfm_3
      + 11'b00000000001;
  assign Gradient_x_calc_COLUMN_acc_5_nl = nl_Gradient_x_calc_COLUMN_acc_5_nl[10:0];
  assign Gradient_x_calc_ROW_not_22_nl = ~ exitL_exit_Gradient_x_calc_ROW_sva;
  assign Gradient_x_calc_ROW_not_21_nl = ~ exitL_exit_Gradient_x_calc_ROW_sva;
  assign Gradient_x_calc_ROW_not_23_nl = ~ exitL_exit_Gradient_x_calc_ROW_sva;
  assign nl_operator_11_false_1_acc_nl = conv_u2u_10_11(Gradient_x_calc_COLUMN_x_lpi_1_dfm_3[10:1])
      + 11'b11111111111;
  assign operator_11_false_1_acc_nl = nl_operator_11_false_1_acc_nl[10:0];
  assign Gradient_x_calc_ROW_not_18_nl = ~ exitL_exit_Gradient_x_calc_ROW_sva;
  assign nl_Gradient_x_calc_COLUMN_acc_8_nl = Gradient_x_calc_COLUMN_mul_itm_1 +
      conv_u2s_34_35({Gradient_x_calc_COLUMN_acc_7_itm_1_33_9 , Gradient_x_calc_COLUMN_acc_7_itm_1_8_0});
  assign Gradient_x_calc_COLUMN_acc_8_nl = nl_Gradient_x_calc_COLUMN_acc_8_nl[34:0];
  assign nl_Gradient_x_calc_COLUMN_acc_9_nl = conv_u2s_37_38(Gradient_x_calc_COLUMN_mul_1_itm_1)
      + conv_s2s_35_38(Gradient_x_calc_COLUMN_acc_8_nl);
  assign Gradient_x_calc_COLUMN_acc_9_nl = nl_Gradient_x_calc_COLUMN_acc_9_nl[37:0];
  assign nl_Gradient_x_calc_COLUMN_acc_nl = Gradient_x_calc_COLUMN_acc_9_nl + Gradient_x_calc_COLUMN_mul_3_itm_1;
  assign Gradient_x_calc_COLUMN_acc_nl = nl_Gradient_x_calc_COLUMN_acc_nl[37:0];
  assign Gradient_x_calc_COLUMN_if_1_not_2_nl = ~ gradient_x_rsci_idat_27_0_mx0c1;

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [27:0] MUX_v_28_2_2;
    input [27:0] input_0;
    input [27:0] input_1;
    input  sel;
    reg [27:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_28_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction


  function automatic [27:0] readslicef_38_28_10;
    input [37:0] vector;
    reg [37:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_38_28_10 = tmp[27:0];
  end
  endfunction


  function automatic [37:0] conv_s2s_35_38 ;
    input [34:0]  vector ;
  begin
    conv_s2s_35_38 = {{3{vector[34]}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [34:0] conv_u2s_34_35 ;
    input [33:0]  vector ;
  begin
    conv_u2s_34_35 =  {1'b0, vector};
  end
  endfunction


  function automatic [37:0] conv_u2s_37_38 ;
    input [36:0]  vector ;
  begin
    conv_u2s_37_38 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_gradient_x_calc
// ------------------------------------------------------------------


module OpticalFlow_gradient_x_calc (
  clk, rst, arst_n, frame3_b_rsc_dat, frame3_b_rsc_vld, frame3_b_rsc_rdy, gradient_x_rsc_dat,
      gradient_x_rsc_vld, gradient_x_rsc_rdy, widthIn, heightIn
);
  input clk;
  input rst;
  input arst_n;
  input [7:0] frame3_b_rsc_dat;
  input frame3_b_rsc_vld;
  output frame3_b_rsc_rdy;
  output [31:0] gradient_x_rsc_dat;
  output gradient_x_rsc_vld;
  input gradient_x_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;



  // Interconnect Declarations for Component Instantiations 
  OpticalFlow_gradient_x_calc_run OpticalFlow_gradient_x_calc_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .frame3_b_rsc_dat(frame3_b_rsc_dat),
      .frame3_b_rsc_vld(frame3_b_rsc_vld),
      .frame3_b_rsc_rdy(frame3_b_rsc_rdy),
      .gradient_x_rsc_dat(gradient_x_rsc_dat),
      .gradient_x_rsc_vld(gradient_x_rsc_vld),
      .gradient_x_rsc_rdy(gradient_x_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn)
    );
endmodule




//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_genreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_genreg_v1 (clk, en, arst, srst, d, z);
    parameter integer width   = 1;
    parameter integer ph_clk  = 1;
    parameter integer ph_en   = 1;
    parameter integer ph_arst = 0;
    parameter integer ph_srst = 1;
    parameter         has_en  = 1'b1;

    input clk;
    input en;
    input arst;
    input srst;
    input      [width-1:0] d;
    output reg [width-1:0] z;

    //  Generate parameters
    //  ph_clk | ph_arst | has_en     Label:
    //    1        1          1       GEN_CLK1_ARST1_EN1
    //    1        1          0       GEN_CLK1_ARST1_EN0
    //    1        0          1       GEN_CLK1_ARST0_EN1
    //    1        0          0       GEN_CLK1_ARST0_EN0
    //    0        1          1       GEN_CLK0_ARST1_EN1
    //    0        1          0       GEN_CLK0_ARST1_EN0
    //    0        0          1       GEN_CLK0_ARST0_EN1
    //    0        0          0       GEN_CLK0_ARST0_EN0
    
    generate 
      // Pos edge clock, pos edge async reset, has enable
      if (ph_clk == 1 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK1_ARST1_EN1
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST1_EN1

      // Pos edge clock, pos edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK1_ARST1_EN0
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST1_EN0

      // Pos edge clock, neg edge async reset, has enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK1_ARST0_EN1
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST0_EN1

      // Pos edge clock, neg edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK1_ARST0_EN0
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST0_EN0


      // Neg edge clock, pos edge async reset, has enable
      if (ph_clk == 0 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK0_ARST1_EN1
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST1_EN1

      // Neg edge clock, pos edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK0_ARST1_EN0
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST1_EN0

      // Neg edge clock, neg edge async reset, has enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK0_ARST0_EN1
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST0_EN1

      // Neg edge clock, neg edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK0_ARST0_EN0
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST0_EN0
    endgenerate
endmodule


//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_fifo_wait_core_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

/*
 *            _________________________________________________
 * WRITER    |                                                 |   READER
 *           |               ccs_fifo_wait_core                |
 *           |             _____________________               |
 *        --<|  din_rdy --<|  ---------------- <|--- dout_rdy <|---
 *           |             |       FIFO         |              |
 *        ---|> din_vld ---|> ----------------  |>-- dout_vld  |>--
 *        ---|>     din ---|> ----------------  |>-- dout      |>--
 *           |             |____________________|              |
 *           |_________________________________________________|
 *
 *    rdy    - can be considered as a notFULL signal
 *    vld    - can be considered as a notEMPTY signal
 *    is_idle - clk can be safely gated
 *
 * Change History:
 *    2019-01-24 - Add assertion to verify rdy signal behavior under reset.
 *                 Fix bug in that behavior.
 */

module ccs_fifo_wait_core_v5 (clk, en, arst, srst, din_vld, din_rdy, din, dout_vld, dout_rdy, dout, sd, is_idle);

    parameter integer rscid    = 0;     // resource ID
    parameter integer width    = 8;     // fifo width
    parameter integer sz_width = 8;     // size of port for elements in fifo
    parameter integer fifo_sz  = 8;     // fifo depth
    parameter integer ph_clk   = 1;     // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1;     // clock enable polarity
    parameter integer ph_arst  = 1;     // async reset polarity
    parameter integer ph_srst  = 1;     // sync reset polarity
    parameter integer ph_log2  = 3;     // log2(fifo_sz)

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 din_vld;    // writer has valid data
    output                din_rdy;    // fifo ready for data (not full)
    input  [width-1:0]    din;
    output                dout_vld;   // fifo has valid data (not empty)
    input                 dout_rdy;   // reader ready for data
    output [width-1:0]    dout;
    output [sz_width-1:0] sd;
    output                is_idle;

    localparam integer fifo_b  = width * fifo_sz;
    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;

    reg      [fifo_mx:0] stat_pre;
    wire     [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [fifo_mx:0] en_l;
    reg      [fifo_mx_over_8:0] en_l_s;

    reg      [width-1:0] buff_nxt;

    reg                  stat_nxt;
    reg                  stat_behind;
    reg                  stat_ahead;
    reg                  stat_tail;
    reg                  en_l_var;

    integer              i;
    genvar               eni;

    wire [32:0]          size_t;
    reg  [31:0]          count;
    reg  [31:0]          count_t;
    reg  [32:0]          n_elem;
    wire                 din_rdy_drv;
    wire                 dout_vld_drv;
    wire                 din_vld_int;
    wire                 hs_init;
    wire                 active;
    wire                 is_idle_drv;

    // synopsys translate_off
    reg  [31:0]          peak;
    initial
    begin
      peak  = 32'b0;
    end
    // synopsys translate_on

    assign din_rdy = din_rdy_drv;
    assign dout_vld = dout_vld_drv;
    assign is_idle = is_idle_drv;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
      assign din_vld_int = din_vld & hs_init;
      assign din_rdy_drv = (dout_rdy | (~stat[0])) & hs_init;
      assign dout_vld_drv = din_vld_int | stat[fifo_sz-1];

      assign active = (din_vld_int & din_rdy_drv) | (dout_rdy & dout_vld_drv);
      assign is_idle_drv = (~active) & hs_init;

      assign size_t = (count - {31'b0, (dout_rdy & stat[fifo_sz-1])}) + {31'b0, din_vld_int};
      assign sd = size_t[sz_width-1:0];

      assign dout = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : din;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_behind = (i != 0) ? stat[i-1] : 1'b0;
          stat_ahead  = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;

          // Determine if this buffer element will have data
          stat_nxt = stat_ahead &                       // valid element ahead of this one (or head)
                       (stat_behind                     // valid element behind this one
                         | (stat[i] & (~dout_rdy))      // valid element and output not ready (in use and not shifted)
                         | (stat[i] & din_vld_int)      // valid element and input has data
                         | (din_vld_int & (~dout_rdy))  // input has data and output not ready
                       );
          stat_pre[i] = stat_nxt;

          // First empty elem when not shifting or last valid elem after shifting (assumes stat_behind == 0)
          stat_tail = stat_ahead & (((~stat[i]) & (~dout_rdy)) | (stat[i] & dout_rdy));

          if (dout_rdy & stat_behind)
          begin
            // shift valid element
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
            en_l_var = 1'b1;
          end
          else if (din_vld_int & stat_tail)
          begin
            // update tail with input data
            buff_nxt = din;
            en_l_var = 1'b1;
          end
          else
          begin
            // no-op, disable register
            buff_nxt = din; // Don't care input to disabled flop
            en_l_var = 1'b0;
          end
          buff_pre[width*i+:width] = buff_nxt[0+:width];

          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          if ((stat_ahead == 1'b1) & (stat[i] == 1'b0))
            //found tail, update the number of elements for count
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end //for loop

        // Enable for stat registers (partitioned into banks of eight)
        // Take care of the head first
        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en & active;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en | ~active;

        // Now every eight
        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if (($unsigned(i) % 32'd8) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]) & (active);
            else
              en_l_s[(i/8)-1] = (en) | (~stat[i]) | (~active);
          end
        end

        // Update count and peak
        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else
          count_t = n_elem[31:0];
        count = count_t;
        // synopsys translate_off
        peak = (peak < count) ? count : peak;
        // synopsys translate_on
      end //FIFOPROC

      // Handshake valid after reset
      ccs_genreg_v1
      #(
        .width   (1),
        .ph_clk  (ph_clk),
        .ph_en   (1),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .has_en  (1'b0)
      )
      HS_INIT_REG
      (
        .clk     (clk),
        .en      (1'b1),
        .arst    (arst),
        .srst    (srst),
        .d       (1'b1),
        .z       (hs_init)
      );

      // Buffer and status registers
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: GEN_REGS
        ccs_genreg_v1
        #(
          .width   (1),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        STATREG
        (
          .clk     (clk),
          .en      (en_l_s[eni/8]),
          .arst    (arst),
          .srst    (srst),
          .d       (stat_pre[eni]),
          .z       (stat[eni])
        );

        ccs_genreg_v1
        #(
          .width   (width),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        BUFREG
        (
          .clk     (clk),
          .en      (en_l[eni]),
          .arst    (arst),
          .srst    (srst),
          .d       (buff_pre[width*eni+:width]),
          .z       (buff[width*eni+:width])
        );
      end

    end
    else
    begin: FEED_THRU
      assign din_rdy_drv  = dout_rdy;
      assign dout_vld_drv = din_vld;
      assign dout     = din;
      // non-blocking is not II=1 when fifo_sz=0
      assign sd = {{(sz_width-1){1'b0}}, (din_vld & ~dout_rdy)};
      assign is_idle_drv = ~(din_vld & dout_rdy);
    end
    endgenerate

`ifdef RDY_ASRT
    generate
    if (ph_clk==1)
    begin: POS_CLK_ASSERT

       property rdyAsrt ;
         @(posedge clk) (srst==ph_srst) |=> (din_rdy==0);
       endproperty
       a1Pos: assert property(rdyAsrt);

       property rdyAsrtASync ;
         @(posedge clk) (arst==ph_arst) |-> (din_rdy==0);
       endproperty
       a2Pos: assert property(rdyAsrtASync);

    end else if (ph_clk==0)
    begin: NEG_CLK_ASSERT

       property rdyAsrt ;
         @(negedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Neg: assert property(rdyAsrt);

       property rdyAsrtASync ;
         @(negedge clk) (arst==ph_arst) |-> (din_rdy==0);
       endproperty
       a2Neg: assert property(rdyAsrtASync);

    end
    endgenerate
`endif

endmodule

//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_pipe_v6.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
/*
 *
 *            _______________________________________________
 * WRITER    |                                              |          READER
 *           |                 ccs_pipe                     |
 *           |            ______________________            |
 *        --<| din_rdy --<|  ---------------- <|---dout_rdy<|---
 *           |            |       FIFO         |            |
 *        ---|>din_vld ---|> ----------------  |>--dout_vld |>--
 *        ---|>din -------|> ----------------  |> -----dout |>--
 *           |            |____________________|            |
 *           |______________________________________________|
 *
 *    din_rdy     - can be considered as a notFULL signal
 *    dout_vld    - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from din_vld & !din_rdy
 *    read_stall  - an internal debug signal formed from dout_rdy & !dout_vld
 *    is_idle     - indicates the clock can be safely gated
 *    stall_ctrl  - Stall the pipe(fifo).  Used by STALL_FLAG_SV directive
 */

module ccs_pipe_v6 (clk, en, arst, srst, din_rdy, din_vld, din, dout_rdy, dout_vld, dout, 
                    sz, sz_req, is_idle);

    parameter integer rscid    = 0; // resource ID
    parameter integer width    = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz  = 8; // fifo depth
    parameter integer log2_sz  = 3; // log2(fifo_sz)
    parameter integer ph_clk   = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1; // clock enable polarity
    parameter integer ph_arst  = 1; // async reset polarity
    parameter integer ph_srst  = 1; // sync reset polarity

    // clock 
    input              clk;
    input              en;
    input              arst;
    input              srst;

    // writer
    output             din_rdy;
    input              din_vld;
    input  [width-1:0] din;

    // reader
    input              dout_rdy;
    output             dout_vld;
    output [width-1:0] dout;

    // size
    output [sz_width-1:0] sz;
    input                 sz_req;
    output                is_idle;

    localparam stallOff = 0; 
    wire                  stall_ctrl;
    assign stall_ctrl = stallOff;
   
    // synopsys translate_off
    wire   write_stall;
    wire   read_stall;
    assign write_stall = (din_vld & !din_rdy) | stall_ctrl;
    assign read_stall  = (dout_rdy & !dout_vld) | stall_ctrl;
    // synopsys translate_on

    wire    tmp_din_rdy;
    assign  din_rdy = tmp_din_rdy & !stall_ctrl;
    wire    tmp_dout_vld;
    assign  dout_vld = tmp_dout_vld & !stall_ctrl;
   
    ccs_fifo_wait_core_v5
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk      (clk),
        .en       (en),
        .arst     (arst),
        .srst     (srst),
        .din_vld  (din_vld & !stall_ctrl),
        .din_rdy  (tmp_din_rdy),
        .din      (din),
        .dout_vld (tmp_dout_vld),
        .dout_rdy (dout_rdy & !stall_ctrl),
        .dout     (dout),
        .sd       (sz),
        .is_idle  (is_idle)
    );

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Mon Jun 17 23:53:59 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    OpticalFlow_Top
// ------------------------------------------------------------------


module OpticalFlow_Top (
  clk, rst, arst_n, input_frames_rsc_dat, input_frames_rsc_vld, input_frames_rsc_rdy,
      widthIn, heightIn, shift_threshold, outputs_rsc_dat, outputs_rsc_vld, outputs_rsc_rdy,
      line_buf3_rsc_clken, line_buf3_rsc_q, line_buf3_rsc_we, line_buf3_rsc_d, line_buf3_rsc_adr,
      line_buf2_rsc_clken, line_buf2_rsc_q, line_buf2_rsc_we, line_buf2_rsc_d, line_buf2_rsc_adr,
      line_buf1_rsc_gradient_y_calc_inst_clken, line_buf1_rsc_gradient_y_calc_inst_q,
      line_buf1_rsc_gradient_y_calc_inst_we, line_buf1_rsc_gradient_y_calc_inst_d,
      line_buf1_rsc_gradient_y_calc_inst_adr, line_buf0_rsc_gradient_y_calc_inst_clken,
      line_buf0_rsc_gradient_y_calc_inst_q, line_buf0_rsc_gradient_y_calc_inst_we,
      line_buf0_rsc_gradient_y_calc_inst_d, line_buf0_rsc_gradient_y_calc_inst_adr,
      line_buf5_Ix_rsc_clken, line_buf5_Ix_rsc_q, line_buf5_Ix_rsc_we, line_buf5_Ix_rsc_d,
      line_buf5_Ix_rsc_adr, line_buf4_Ix_rsc_clken, line_buf4_Ix_rsc_q, line_buf4_Ix_rsc_we,
      line_buf4_Ix_rsc_d, line_buf4_Ix_rsc_adr, line_buf3_Ix_rsc_clken, line_buf3_Ix_rsc_q,
      line_buf3_Ix_rsc_we, line_buf3_Ix_rsc_d, line_buf3_Ix_rsc_adr, line_buf2_Ix_rsc_clken,
      line_buf2_Ix_rsc_q, line_buf2_Ix_rsc_we, line_buf2_Ix_rsc_d, line_buf2_Ix_rsc_adr,
      line_buf1_Ix_rsc_clken, line_buf1_Ix_rsc_q, line_buf1_Ix_rsc_we, line_buf1_Ix_rsc_d,
      line_buf1_Ix_rsc_adr, line_buf0_Ix_rsc_clken, line_buf0_Ix_rsc_q, line_buf0_Ix_rsc_we,
      line_buf0_Ix_rsc_d, line_buf0_Ix_rsc_adr, line_buf5_Iy_rsc_clken, line_buf5_Iy_rsc_q,
      line_buf5_Iy_rsc_we, line_buf5_Iy_rsc_d, line_buf5_Iy_rsc_adr, line_buf4_Iy_rsc_clken,
      line_buf4_Iy_rsc_q, line_buf4_Iy_rsc_we, line_buf4_Iy_rsc_d, line_buf4_Iy_rsc_adr,
      line_buf3_Iy_rsc_clken, line_buf3_Iy_rsc_q, line_buf3_Iy_rsc_we, line_buf3_Iy_rsc_d,
      line_buf3_Iy_rsc_adr, line_buf2_Iy_rsc_clken, line_buf2_Iy_rsc_q, line_buf2_Iy_rsc_we,
      line_buf2_Iy_rsc_d, line_buf2_Iy_rsc_adr, line_buf1_Iy_rsc_clken, line_buf1_Iy_rsc_q,
      line_buf1_Iy_rsc_we, line_buf1_Iy_rsc_d, line_buf1_Iy_rsc_adr, line_buf0_Iy_rsc_clken,
      line_buf0_Iy_rsc_q, line_buf0_Iy_rsc_we, line_buf0_Iy_rsc_d, line_buf0_Iy_rsc_adr,
      line_buf5_Iz_rsc_clken, line_buf5_Iz_rsc_q, line_buf5_Iz_rsc_we, line_buf5_Iz_rsc_d,
      line_buf5_Iz_rsc_adr, line_buf4_Iz_rsc_clken, line_buf4_Iz_rsc_q, line_buf4_Iz_rsc_we,
      line_buf4_Iz_rsc_d, line_buf4_Iz_rsc_adr, line_buf3_Iz_rsc_clken, line_buf3_Iz_rsc_q,
      line_buf3_Iz_rsc_we, line_buf3_Iz_rsc_d, line_buf3_Iz_rsc_adr, line_buf2_Iz_rsc_clken,
      line_buf2_Iz_rsc_q, line_buf2_Iz_rsc_we, line_buf2_Iz_rsc_d, line_buf2_Iz_rsc_adr,
      line_buf1_Iz_rsc_clken, line_buf1_Iz_rsc_q, line_buf1_Iz_rsc_we, line_buf1_Iz_rsc_d,
      line_buf1_Iz_rsc_adr, line_buf0_Iz_rsc_clken, line_buf0_Iz_rsc_q, line_buf0_Iz_rsc_we,
      line_buf0_Iz_rsc_d, line_buf0_Iz_rsc_adr, line_buf1_rsc_tensor_weight_y_inst_clken,
      line_buf1_rsc_tensor_weight_y_inst_q, line_buf1_rsc_tensor_weight_y_inst_we,
      line_buf1_rsc_tensor_weight_y_inst_d, line_buf1_rsc_tensor_weight_y_inst_adr,
      line_buf0_rsc_tensor_weight_y_inst_clken, line_buf0_rsc_tensor_weight_y_inst_q,
      line_buf0_rsc_tensor_weight_y_inst_we, line_buf0_rsc_tensor_weight_y_inst_d,
      line_buf0_rsc_tensor_weight_y_inst_adr
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] input_frames_rsc_dat;
  input input_frames_rsc_vld;
  output input_frames_rsc_rdy;
  input [10:0] widthIn;
  input [8:0] heightIn;
  input [8:0] shift_threshold;
  output [31:0] outputs_rsc_dat;
  output outputs_rsc_vld;
  input outputs_rsc_rdy;
  output line_buf3_rsc_clken;
  input [15:0] line_buf3_rsc_q;
  output line_buf3_rsc_we;
  output [15:0] line_buf3_rsc_d;
  output [8:0] line_buf3_rsc_adr;
  output line_buf2_rsc_clken;
  input [15:0] line_buf2_rsc_q;
  output line_buf2_rsc_we;
  output [15:0] line_buf2_rsc_d;
  output [8:0] line_buf2_rsc_adr;
  output line_buf1_rsc_gradient_y_calc_inst_clken;
  input [63:0] line_buf1_rsc_gradient_y_calc_inst_q;
  output line_buf1_rsc_gradient_y_calc_inst_we;
  output [63:0] line_buf1_rsc_gradient_y_calc_inst_d;
  output [8:0] line_buf1_rsc_gradient_y_calc_inst_adr;
  output line_buf0_rsc_gradient_y_calc_inst_clken;
  input [63:0] line_buf0_rsc_gradient_y_calc_inst_q;
  output line_buf0_rsc_gradient_y_calc_inst_we;
  output [63:0] line_buf0_rsc_gradient_y_calc_inst_d;
  output [8:0] line_buf0_rsc_gradient_y_calc_inst_adr;
  output line_buf5_Ix_rsc_clken;
  input [63:0] line_buf5_Ix_rsc_q;
  output line_buf5_Ix_rsc_we;
  output [63:0] line_buf5_Ix_rsc_d;
  output [8:0] line_buf5_Ix_rsc_adr;
  output line_buf4_Ix_rsc_clken;
  input [63:0] line_buf4_Ix_rsc_q;
  output line_buf4_Ix_rsc_we;
  output [63:0] line_buf4_Ix_rsc_d;
  output [8:0] line_buf4_Ix_rsc_adr;
  output line_buf3_Ix_rsc_clken;
  input [63:0] line_buf3_Ix_rsc_q;
  output line_buf3_Ix_rsc_we;
  output [63:0] line_buf3_Ix_rsc_d;
  output [8:0] line_buf3_Ix_rsc_adr;
  output line_buf2_Ix_rsc_clken;
  input [63:0] line_buf2_Ix_rsc_q;
  output line_buf2_Ix_rsc_we;
  output [63:0] line_buf2_Ix_rsc_d;
  output [8:0] line_buf2_Ix_rsc_adr;
  output line_buf1_Ix_rsc_clken;
  input [63:0] line_buf1_Ix_rsc_q;
  output line_buf1_Ix_rsc_we;
  output [63:0] line_buf1_Ix_rsc_d;
  output [8:0] line_buf1_Ix_rsc_adr;
  output line_buf0_Ix_rsc_clken;
  input [63:0] line_buf0_Ix_rsc_q;
  output line_buf0_Ix_rsc_we;
  output [63:0] line_buf0_Ix_rsc_d;
  output [8:0] line_buf0_Ix_rsc_adr;
  output line_buf5_Iy_rsc_clken;
  input [63:0] line_buf5_Iy_rsc_q;
  output line_buf5_Iy_rsc_we;
  output [63:0] line_buf5_Iy_rsc_d;
  output [8:0] line_buf5_Iy_rsc_adr;
  output line_buf4_Iy_rsc_clken;
  input [63:0] line_buf4_Iy_rsc_q;
  output line_buf4_Iy_rsc_we;
  output [63:0] line_buf4_Iy_rsc_d;
  output [8:0] line_buf4_Iy_rsc_adr;
  output line_buf3_Iy_rsc_clken;
  input [63:0] line_buf3_Iy_rsc_q;
  output line_buf3_Iy_rsc_we;
  output [63:0] line_buf3_Iy_rsc_d;
  output [8:0] line_buf3_Iy_rsc_adr;
  output line_buf2_Iy_rsc_clken;
  input [63:0] line_buf2_Iy_rsc_q;
  output line_buf2_Iy_rsc_we;
  output [63:0] line_buf2_Iy_rsc_d;
  output [8:0] line_buf2_Iy_rsc_adr;
  output line_buf1_Iy_rsc_clken;
  input [63:0] line_buf1_Iy_rsc_q;
  output line_buf1_Iy_rsc_we;
  output [63:0] line_buf1_Iy_rsc_d;
  output [8:0] line_buf1_Iy_rsc_adr;
  output line_buf0_Iy_rsc_clken;
  input [63:0] line_buf0_Iy_rsc_q;
  output line_buf0_Iy_rsc_we;
  output [63:0] line_buf0_Iy_rsc_d;
  output [8:0] line_buf0_Iy_rsc_adr;
  output line_buf5_Iz_rsc_clken;
  input [63:0] line_buf5_Iz_rsc_q;
  output line_buf5_Iz_rsc_we;
  output [63:0] line_buf5_Iz_rsc_d;
  output [8:0] line_buf5_Iz_rsc_adr;
  output line_buf4_Iz_rsc_clken;
  input [63:0] line_buf4_Iz_rsc_q;
  output line_buf4_Iz_rsc_we;
  output [63:0] line_buf4_Iz_rsc_d;
  output [8:0] line_buf4_Iz_rsc_adr;
  output line_buf3_Iz_rsc_clken;
  input [63:0] line_buf3_Iz_rsc_q;
  output line_buf3_Iz_rsc_we;
  output [63:0] line_buf3_Iz_rsc_d;
  output [8:0] line_buf3_Iz_rsc_adr;
  output line_buf2_Iz_rsc_clken;
  input [63:0] line_buf2_Iz_rsc_q;
  output line_buf2_Iz_rsc_we;
  output [63:0] line_buf2_Iz_rsc_d;
  output [8:0] line_buf2_Iz_rsc_adr;
  output line_buf1_Iz_rsc_clken;
  input [63:0] line_buf1_Iz_rsc_q;
  output line_buf1_Iz_rsc_we;
  output [63:0] line_buf1_Iz_rsc_d;
  output [8:0] line_buf1_Iz_rsc_adr;
  output line_buf0_Iz_rsc_clken;
  input [63:0] line_buf0_Iz_rsc_q;
  output line_buf0_Iz_rsc_we;
  output [63:0] line_buf0_Iz_rsc_d;
  output [8:0] line_buf0_Iz_rsc_adr;
  output line_buf1_rsc_tensor_weight_y_inst_clken;
  input [767:0] line_buf1_rsc_tensor_weight_y_inst_q;
  output line_buf1_rsc_tensor_weight_y_inst_we;
  output [767:0] line_buf1_rsc_tensor_weight_y_inst_d;
  output [8:0] line_buf1_rsc_tensor_weight_y_inst_adr;
  output line_buf0_rsc_tensor_weight_y_inst_clken;
  input [767:0] line_buf0_rsc_tensor_weight_y_inst_q;
  output line_buf0_rsc_tensor_weight_y_inst_we;
  output [767:0] line_buf0_rsc_tensor_weight_y_inst_d;
  output [8:0] line_buf0_rsc_tensor_weight_y_inst_adr;


  // Interconnect Declarations
  wire [31:0] gradient_x_rsc_dat_n_gradient_x_calc_inst;
  wire [31:0] gradient_y_rsc_dat_n_gradient_y_calc_inst;
  wire gradient_y_rsc_rdy_n_gradient_y_calc_inst;
  wire [7:0] frame3_rsc_dat_n_gradient_y_calc_inst;
  wire [31:0] input_frames_delayed_rsc_dat_n_gradient_y_calc_inst;
  wire line_buf3_rsc_clken_n_gradient_y_calc_inst;
  wire [15:0] line_buf3_rsc_d_n_gradient_y_calc_inst;
  wire [8:0] line_buf3_rsc_adr_n_gradient_y_calc_inst;
  wire line_buf2_rsc_clken_n_gradient_y_calc_inst;
  wire [15:0] line_buf2_rsc_d_n_gradient_y_calc_inst;
  wire [8:0] line_buf2_rsc_adr_n_gradient_y_calc_inst;
  wire line_buf1_rsc_clken_n_gradient_y_calc_inst;
  wire [63:0] line_buf1_rsc_d_n_gradient_y_calc_inst;
  wire [8:0] line_buf1_rsc_adr_n_gradient_y_calc_inst;
  wire line_buf0_rsc_clken_n_gradient_y_calc_inst;
  wire [63:0] line_buf0_rsc_d_n_gradient_y_calc_inst;
  wire [8:0] line_buf0_rsc_adr_n_gradient_y_calc_inst;
  wire [31:0] gradient_z_rsc_dat_n_gradient_z_calc_inst;
  wire gradient_z_rsc_rdy_n_gradient_z_calc_inst;
  wire [31:0] gradient_y_rsc_dat_n_gradient_weight_y_inst;
  wire gradient_y_rsc_vld_n_gradient_weight_y_inst;
  wire [31:0] gradient_z_rsc_dat_n_gradient_weight_y_inst;
  wire gradient_z_rsc_vld_n_gradient_weight_y_inst;
  wire [95:0] y_filtered_rsc_dat_n_gradient_weight_y_inst;
  wire line_buf5_Ix_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf5_Ix_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf5_Ix_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf4_Ix_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf4_Ix_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf4_Ix_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf3_Ix_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf3_Ix_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf3_Ix_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf2_Ix_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf2_Ix_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf2_Ix_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf1_Ix_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf1_Ix_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf1_Ix_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf0_Ix_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf0_Ix_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf0_Ix_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf5_Iy_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf5_Iy_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf5_Iy_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf4_Iy_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf4_Iy_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf4_Iy_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf3_Iy_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf3_Iy_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf3_Iy_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf2_Iy_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf2_Iy_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf2_Iy_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf1_Iy_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf1_Iy_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf1_Iy_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf0_Iy_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf0_Iy_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf0_Iy_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf5_Iz_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf5_Iz_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf5_Iz_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf4_Iz_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf4_Iz_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf4_Iz_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf3_Iz_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf3_Iz_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf3_Iz_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf2_Iz_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf2_Iz_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf2_Iz_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf1_Iz_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf1_Iz_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf1_Iz_rsc_adr_n_gradient_weight_y_inst;
  wire line_buf0_Iz_rsc_clken_n_gradient_weight_y_inst;
  wire [63:0] line_buf0_Iz_rsc_d_n_gradient_weight_y_inst;
  wire [8:0] line_buf0_Iz_rsc_adr_n_gradient_weight_y_inst;
  wire [95:0] filtered_gradient_rsc_dat_n_gradient_weight_x_inst;
  wire [383:0] out_product_rsc_dat_n_outer_product_inst;
  wire [383:0] tensor_y_rsc_dat_n_tensor_weight_y_inst;
  wire line_buf1_rsc_clken_n_tensor_weight_y_inst;
  wire [767:0] line_buf1_rsc_d_n_tensor_weight_y_inst;
  wire [8:0] line_buf1_rsc_adr_n_tensor_weight_y_inst;
  wire line_buf0_rsc_clken_n_tensor_weight_y_inst;
  wire [767:0] line_buf0_rsc_d_n_tensor_weight_y_inst;
  wire [8:0] line_buf0_rsc_adr_n_tensor_weight_y_inst;
  wire [191:0] tensor_shift_rsc_dat_n_tensor_weight_x_inst;
  wire [8:0] shift_rsc_dat_n_tensor_weight_x_inst;
  wire [31:0] output_rsc_dat_n_flow_calc_inst;
  wire frame3_b_rsc_rdy_n_gradient_x_calc_inst_bud;
  wire frame3_rsc_vld_n_gradient_y_calc_inst_bud;
  wire gradient_x_rsc_vld_n_gradient_x_calc_inst_bud;
  wire gradient_x_rsc_rdy_n_gradient_weight_y_inst_bud;
  wire input_frames_rsc_rdy_n_gradient_y_calc_inst_bud;
  wire gradient_y_rsc_vld_n_gradient_y_calc_inst_bud;
  wire gradient_y_rsc_rdy_n_gradient_weight_y_inst_bud;
  wire input_frames_delayed_rsc_vld_n_gradient_y_calc_inst_bud;
  wire input_frames_delayed_rsc_rdy_n_gradient_z_calc_inst_bud;
  wire line_buf3_rsc_we_n_gradient_y_calc_inst_bud;
  wire line_buf2_rsc_we_n_gradient_y_calc_inst_bud;
  wire line_buf1_rsc_we_n_gradient_y_calc_inst_bud;
  wire line_buf0_rsc_we_n_gradient_y_calc_inst_bud;
  wire gradient_z_rsc_vld_n_gradient_z_calc_inst_bud;
  wire gradient_z_rsc_rdy_n_gradient_weight_y_inst_bud;
  wire y_filtered_rsc_vld_n_gradient_weight_y_inst_bud;
  wire y_filtered_rsc_rdy_n_gradient_weight_x_inst_bud;
  wire line_buf5_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf4_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf3_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf2_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf1_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf0_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf5_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf4_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf3_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf2_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf1_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf0_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf5_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf4_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf3_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf2_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf1_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  wire line_buf0_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  wire filtered_gradient_rsc_vld_n_gradient_weight_x_inst_bud;
  wire filtered_gradient_rsc_rdy_n_outer_product_inst_bud;
  wire out_product_rsc_vld_n_outer_product_inst_bud;
  wire out_product_rsc_rdy_n_tensor_weight_y_inst_bud;
  wire tensor_y_rsc_vld_n_tensor_weight_y_inst_bud;
  wire tensor_y_rsc_rdy_n_tensor_weight_x_inst_bud;
  wire line_buf1_rsc_we_n_tensor_weight_y_inst_bud;
  wire line_buf0_rsc_we_n_tensor_weight_y_inst_bud;
  wire tensor_shift_rsc_vld_n_tensor_weight_x_inst_bud;
  wire tensor_shift_rsc_rdy_n_flow_calc_inst_bud;
  wire shift_rsc_vld_n_tensor_weight_x_inst_bud;
  wire shift_rsc_rdy_n_flow_calc_inst_bud;
  wire output_rsc_vld_n_flow_calc_inst_bud;
  wire gradient_y_unc_1;
  wire gradient_y_idle;
  wire gradient_z_unc_1;
  wire gradient_z_idle;


  // Interconnect Declarations for Component Instantiations 
  ccs_pipe_v6 #(.rscid(32'sd87),
  .width(32'sd32),
  .sz_width(32'sd1),
  .fifo_sz(32'sd4),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd1)) gradient_y_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(rst),
      .din_rdy(gradient_y_rsc_rdy_n_gradient_y_calc_inst),
      .din_vld(gradient_y_rsc_vld_n_gradient_y_calc_inst_bud),
      .din(gradient_y_rsc_dat_n_gradient_y_calc_inst),
      .dout_rdy(gradient_y_rsc_rdy_n_gradient_weight_y_inst_bud),
      .dout_vld(gradient_y_rsc_vld_n_gradient_weight_y_inst),
      .dout(gradient_y_rsc_dat_n_gradient_weight_y_inst),
      .sz(gradient_y_unc_1),
      .sz_req(1'b0),
      .is_idle(gradient_y_idle)
    );
  ccs_pipe_v6 #(.rscid(32'sd88),
  .width(32'sd32),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd1)) gradient_z_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(rst),
      .din_rdy(gradient_z_rsc_rdy_n_gradient_z_calc_inst),
      .din_vld(gradient_z_rsc_vld_n_gradient_z_calc_inst_bud),
      .din(gradient_z_rsc_dat_n_gradient_z_calc_inst),
      .dout_rdy(gradient_z_rsc_rdy_n_gradient_weight_y_inst_bud),
      .dout_vld(gradient_z_rsc_vld_n_gradient_weight_y_inst),
      .dout(gradient_z_rsc_dat_n_gradient_weight_y_inst),
      .sz(gradient_z_unc_1),
      .sz_req(1'b0),
      .is_idle(gradient_z_idle)
    );
  OpticalFlow_gradient_x_calc gradient_x_calc_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .frame3_b_rsc_dat(frame3_rsc_dat_n_gradient_y_calc_inst),
      .frame3_b_rsc_vld(frame3_rsc_vld_n_gradient_y_calc_inst_bud),
      .frame3_b_rsc_rdy(frame3_b_rsc_rdy_n_gradient_x_calc_inst_bud),
      .gradient_x_rsc_dat(gradient_x_rsc_dat_n_gradient_x_calc_inst),
      .gradient_x_rsc_vld(gradient_x_rsc_vld_n_gradient_x_calc_inst_bud),
      .gradient_x_rsc_rdy(gradient_x_rsc_rdy_n_gradient_weight_y_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn)
    );
  OpticalFlow_gradient_y_calc gradient_y_calc_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .input_frames_rsc_dat(input_frames_rsc_dat),
      .input_frames_rsc_vld(input_frames_rsc_vld),
      .input_frames_rsc_rdy(input_frames_rsc_rdy_n_gradient_y_calc_inst_bud),
      .gradient_y_rsc_dat(gradient_y_rsc_dat_n_gradient_y_calc_inst),
      .gradient_y_rsc_vld(gradient_y_rsc_vld_n_gradient_y_calc_inst_bud),
      .gradient_y_rsc_rdy(gradient_y_rsc_rdy_n_gradient_y_calc_inst),
      .frame3_rsc_dat(frame3_rsc_dat_n_gradient_y_calc_inst),
      .frame3_rsc_vld(frame3_rsc_vld_n_gradient_y_calc_inst_bud),
      .frame3_rsc_rdy(frame3_b_rsc_rdy_n_gradient_x_calc_inst_bud),
      .input_frames_delayed_rsc_dat(input_frames_delayed_rsc_dat_n_gradient_y_calc_inst),
      .input_frames_delayed_rsc_vld(input_frames_delayed_rsc_vld_n_gradient_y_calc_inst_bud),
      .input_frames_delayed_rsc_rdy(input_frames_delayed_rsc_rdy_n_gradient_z_calc_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .line_buf3_rsc_clken(line_buf3_rsc_clken_n_gradient_y_calc_inst),
      .line_buf3_rsc_q(line_buf3_rsc_q),
      .line_buf3_rsc_we(line_buf3_rsc_we_n_gradient_y_calc_inst_bud),
      .line_buf3_rsc_d(line_buf3_rsc_d_n_gradient_y_calc_inst),
      .line_buf3_rsc_adr(line_buf3_rsc_adr_n_gradient_y_calc_inst),
      .line_buf2_rsc_clken(line_buf2_rsc_clken_n_gradient_y_calc_inst),
      .line_buf2_rsc_q(line_buf2_rsc_q),
      .line_buf2_rsc_we(line_buf2_rsc_we_n_gradient_y_calc_inst_bud),
      .line_buf2_rsc_d(line_buf2_rsc_d_n_gradient_y_calc_inst),
      .line_buf2_rsc_adr(line_buf2_rsc_adr_n_gradient_y_calc_inst),
      .line_buf1_rsc_clken(line_buf1_rsc_clken_n_gradient_y_calc_inst),
      .line_buf1_rsc_q(line_buf1_rsc_gradient_y_calc_inst_q),
      .line_buf1_rsc_we(line_buf1_rsc_we_n_gradient_y_calc_inst_bud),
      .line_buf1_rsc_d(line_buf1_rsc_d_n_gradient_y_calc_inst),
      .line_buf1_rsc_adr(line_buf1_rsc_adr_n_gradient_y_calc_inst),
      .line_buf0_rsc_clken(line_buf0_rsc_clken_n_gradient_y_calc_inst),
      .line_buf0_rsc_q(line_buf0_rsc_gradient_y_calc_inst_q),
      .line_buf0_rsc_we(line_buf0_rsc_we_n_gradient_y_calc_inst_bud),
      .line_buf0_rsc_d(line_buf0_rsc_d_n_gradient_y_calc_inst),
      .line_buf0_rsc_adr(line_buf0_rsc_adr_n_gradient_y_calc_inst)
    );
  OpticalFlow_gradient_z_calc gradient_z_calc_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .input_frames_delayed_rsc_dat(input_frames_delayed_rsc_dat_n_gradient_y_calc_inst),
      .input_frames_delayed_rsc_vld(input_frames_delayed_rsc_vld_n_gradient_y_calc_inst_bud),
      .input_frames_delayed_rsc_rdy(input_frames_delayed_rsc_rdy_n_gradient_z_calc_inst_bud),
      .gradient_z_rsc_dat(gradient_z_rsc_dat_n_gradient_z_calc_inst),
      .gradient_z_rsc_vld(gradient_z_rsc_vld_n_gradient_z_calc_inst_bud),
      .gradient_z_rsc_rdy(gradient_z_rsc_rdy_n_gradient_z_calc_inst),
      .widthIn(widthIn),
      .heightIn(heightIn)
    );
  OpticalFlow_gradient_weight_y gradient_weight_y_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .gradient_x_rsc_dat(gradient_x_rsc_dat_n_gradient_x_calc_inst),
      .gradient_x_rsc_vld(gradient_x_rsc_vld_n_gradient_x_calc_inst_bud),
      .gradient_x_rsc_rdy(gradient_x_rsc_rdy_n_gradient_weight_y_inst_bud),
      .gradient_y_rsc_dat(gradient_y_rsc_dat_n_gradient_weight_y_inst),
      .gradient_y_rsc_vld(gradient_y_rsc_vld_n_gradient_weight_y_inst),
      .gradient_y_rsc_rdy(gradient_y_rsc_rdy_n_gradient_weight_y_inst_bud),
      .gradient_z_rsc_dat(gradient_z_rsc_dat_n_gradient_weight_y_inst),
      .gradient_z_rsc_vld(gradient_z_rsc_vld_n_gradient_weight_y_inst),
      .gradient_z_rsc_rdy(gradient_z_rsc_rdy_n_gradient_weight_y_inst_bud),
      .y_filtered_rsc_dat(y_filtered_rsc_dat_n_gradient_weight_y_inst),
      .y_filtered_rsc_vld(y_filtered_rsc_vld_n_gradient_weight_y_inst_bud),
      .y_filtered_rsc_rdy(y_filtered_rsc_rdy_n_gradient_weight_x_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .line_buf5_Ix_rsc_clken(line_buf5_Ix_rsc_clken_n_gradient_weight_y_inst),
      .line_buf5_Ix_rsc_q(line_buf5_Ix_rsc_q),
      .line_buf5_Ix_rsc_we(line_buf5_Ix_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf5_Ix_rsc_d(line_buf5_Ix_rsc_d_n_gradient_weight_y_inst),
      .line_buf5_Ix_rsc_adr(line_buf5_Ix_rsc_adr_n_gradient_weight_y_inst),
      .line_buf4_Ix_rsc_clken(line_buf4_Ix_rsc_clken_n_gradient_weight_y_inst),
      .line_buf4_Ix_rsc_q(line_buf4_Ix_rsc_q),
      .line_buf4_Ix_rsc_we(line_buf4_Ix_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf4_Ix_rsc_d(line_buf4_Ix_rsc_d_n_gradient_weight_y_inst),
      .line_buf4_Ix_rsc_adr(line_buf4_Ix_rsc_adr_n_gradient_weight_y_inst),
      .line_buf3_Ix_rsc_clken(line_buf3_Ix_rsc_clken_n_gradient_weight_y_inst),
      .line_buf3_Ix_rsc_q(line_buf3_Ix_rsc_q),
      .line_buf3_Ix_rsc_we(line_buf3_Ix_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf3_Ix_rsc_d(line_buf3_Ix_rsc_d_n_gradient_weight_y_inst),
      .line_buf3_Ix_rsc_adr(line_buf3_Ix_rsc_adr_n_gradient_weight_y_inst),
      .line_buf2_Ix_rsc_clken(line_buf2_Ix_rsc_clken_n_gradient_weight_y_inst),
      .line_buf2_Ix_rsc_q(line_buf2_Ix_rsc_q),
      .line_buf2_Ix_rsc_we(line_buf2_Ix_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf2_Ix_rsc_d(line_buf2_Ix_rsc_d_n_gradient_weight_y_inst),
      .line_buf2_Ix_rsc_adr(line_buf2_Ix_rsc_adr_n_gradient_weight_y_inst),
      .line_buf1_Ix_rsc_clken(line_buf1_Ix_rsc_clken_n_gradient_weight_y_inst),
      .line_buf1_Ix_rsc_q(line_buf1_Ix_rsc_q),
      .line_buf1_Ix_rsc_we(line_buf1_Ix_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf1_Ix_rsc_d(line_buf1_Ix_rsc_d_n_gradient_weight_y_inst),
      .line_buf1_Ix_rsc_adr(line_buf1_Ix_rsc_adr_n_gradient_weight_y_inst),
      .line_buf0_Ix_rsc_clken(line_buf0_Ix_rsc_clken_n_gradient_weight_y_inst),
      .line_buf0_Ix_rsc_q(line_buf0_Ix_rsc_q),
      .line_buf0_Ix_rsc_we(line_buf0_Ix_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf0_Ix_rsc_d(line_buf0_Ix_rsc_d_n_gradient_weight_y_inst),
      .line_buf0_Ix_rsc_adr(line_buf0_Ix_rsc_adr_n_gradient_weight_y_inst),
      .line_buf5_Iy_rsc_clken(line_buf5_Iy_rsc_clken_n_gradient_weight_y_inst),
      .line_buf5_Iy_rsc_q(line_buf5_Iy_rsc_q),
      .line_buf5_Iy_rsc_we(line_buf5_Iy_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf5_Iy_rsc_d(line_buf5_Iy_rsc_d_n_gradient_weight_y_inst),
      .line_buf5_Iy_rsc_adr(line_buf5_Iy_rsc_adr_n_gradient_weight_y_inst),
      .line_buf4_Iy_rsc_clken(line_buf4_Iy_rsc_clken_n_gradient_weight_y_inst),
      .line_buf4_Iy_rsc_q(line_buf4_Iy_rsc_q),
      .line_buf4_Iy_rsc_we(line_buf4_Iy_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf4_Iy_rsc_d(line_buf4_Iy_rsc_d_n_gradient_weight_y_inst),
      .line_buf4_Iy_rsc_adr(line_buf4_Iy_rsc_adr_n_gradient_weight_y_inst),
      .line_buf3_Iy_rsc_clken(line_buf3_Iy_rsc_clken_n_gradient_weight_y_inst),
      .line_buf3_Iy_rsc_q(line_buf3_Iy_rsc_q),
      .line_buf3_Iy_rsc_we(line_buf3_Iy_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf3_Iy_rsc_d(line_buf3_Iy_rsc_d_n_gradient_weight_y_inst),
      .line_buf3_Iy_rsc_adr(line_buf3_Iy_rsc_adr_n_gradient_weight_y_inst),
      .line_buf2_Iy_rsc_clken(line_buf2_Iy_rsc_clken_n_gradient_weight_y_inst),
      .line_buf2_Iy_rsc_q(line_buf2_Iy_rsc_q),
      .line_buf2_Iy_rsc_we(line_buf2_Iy_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf2_Iy_rsc_d(line_buf2_Iy_rsc_d_n_gradient_weight_y_inst),
      .line_buf2_Iy_rsc_adr(line_buf2_Iy_rsc_adr_n_gradient_weight_y_inst),
      .line_buf1_Iy_rsc_clken(line_buf1_Iy_rsc_clken_n_gradient_weight_y_inst),
      .line_buf1_Iy_rsc_q(line_buf1_Iy_rsc_q),
      .line_buf1_Iy_rsc_we(line_buf1_Iy_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf1_Iy_rsc_d(line_buf1_Iy_rsc_d_n_gradient_weight_y_inst),
      .line_buf1_Iy_rsc_adr(line_buf1_Iy_rsc_adr_n_gradient_weight_y_inst),
      .line_buf0_Iy_rsc_clken(line_buf0_Iy_rsc_clken_n_gradient_weight_y_inst),
      .line_buf0_Iy_rsc_q(line_buf0_Iy_rsc_q),
      .line_buf0_Iy_rsc_we(line_buf0_Iy_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf0_Iy_rsc_d(line_buf0_Iy_rsc_d_n_gradient_weight_y_inst),
      .line_buf0_Iy_rsc_adr(line_buf0_Iy_rsc_adr_n_gradient_weight_y_inst),
      .line_buf5_Iz_rsc_clken(line_buf5_Iz_rsc_clken_n_gradient_weight_y_inst),
      .line_buf5_Iz_rsc_q(line_buf5_Iz_rsc_q),
      .line_buf5_Iz_rsc_we(line_buf5_Iz_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf5_Iz_rsc_d(line_buf5_Iz_rsc_d_n_gradient_weight_y_inst),
      .line_buf5_Iz_rsc_adr(line_buf5_Iz_rsc_adr_n_gradient_weight_y_inst),
      .line_buf4_Iz_rsc_clken(line_buf4_Iz_rsc_clken_n_gradient_weight_y_inst),
      .line_buf4_Iz_rsc_q(line_buf4_Iz_rsc_q),
      .line_buf4_Iz_rsc_we(line_buf4_Iz_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf4_Iz_rsc_d(line_buf4_Iz_rsc_d_n_gradient_weight_y_inst),
      .line_buf4_Iz_rsc_adr(line_buf4_Iz_rsc_adr_n_gradient_weight_y_inst),
      .line_buf3_Iz_rsc_clken(line_buf3_Iz_rsc_clken_n_gradient_weight_y_inst),
      .line_buf3_Iz_rsc_q(line_buf3_Iz_rsc_q),
      .line_buf3_Iz_rsc_we(line_buf3_Iz_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf3_Iz_rsc_d(line_buf3_Iz_rsc_d_n_gradient_weight_y_inst),
      .line_buf3_Iz_rsc_adr(line_buf3_Iz_rsc_adr_n_gradient_weight_y_inst),
      .line_buf2_Iz_rsc_clken(line_buf2_Iz_rsc_clken_n_gradient_weight_y_inst),
      .line_buf2_Iz_rsc_q(line_buf2_Iz_rsc_q),
      .line_buf2_Iz_rsc_we(line_buf2_Iz_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf2_Iz_rsc_d(line_buf2_Iz_rsc_d_n_gradient_weight_y_inst),
      .line_buf2_Iz_rsc_adr(line_buf2_Iz_rsc_adr_n_gradient_weight_y_inst),
      .line_buf1_Iz_rsc_clken(line_buf1_Iz_rsc_clken_n_gradient_weight_y_inst),
      .line_buf1_Iz_rsc_q(line_buf1_Iz_rsc_q),
      .line_buf1_Iz_rsc_we(line_buf1_Iz_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf1_Iz_rsc_d(line_buf1_Iz_rsc_d_n_gradient_weight_y_inst),
      .line_buf1_Iz_rsc_adr(line_buf1_Iz_rsc_adr_n_gradient_weight_y_inst),
      .line_buf0_Iz_rsc_clken(line_buf0_Iz_rsc_clken_n_gradient_weight_y_inst),
      .line_buf0_Iz_rsc_q(line_buf0_Iz_rsc_q),
      .line_buf0_Iz_rsc_we(line_buf0_Iz_rsc_we_n_gradient_weight_y_inst_bud),
      .line_buf0_Iz_rsc_d(line_buf0_Iz_rsc_d_n_gradient_weight_y_inst),
      .line_buf0_Iz_rsc_adr(line_buf0_Iz_rsc_adr_n_gradient_weight_y_inst)
    );
  OpticalFlow_gradient_weight_x gradient_weight_x_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .y_filtered_rsc_dat(y_filtered_rsc_dat_n_gradient_weight_y_inst),
      .y_filtered_rsc_vld(y_filtered_rsc_vld_n_gradient_weight_y_inst_bud),
      .y_filtered_rsc_rdy(y_filtered_rsc_rdy_n_gradient_weight_x_inst_bud),
      .filtered_gradient_rsc_dat(filtered_gradient_rsc_dat_n_gradient_weight_x_inst),
      .filtered_gradient_rsc_vld(filtered_gradient_rsc_vld_n_gradient_weight_x_inst_bud),
      .filtered_gradient_rsc_rdy(filtered_gradient_rsc_rdy_n_outer_product_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn)
    );
  OpticalFlow_outer_product outer_product_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .filtered_gradient_rsc_dat(filtered_gradient_rsc_dat_n_gradient_weight_x_inst),
      .filtered_gradient_rsc_vld(filtered_gradient_rsc_vld_n_gradient_weight_x_inst_bud),
      .filtered_gradient_rsc_rdy(filtered_gradient_rsc_rdy_n_outer_product_inst_bud),
      .out_product_rsc_dat(out_product_rsc_dat_n_outer_product_inst),
      .out_product_rsc_vld(out_product_rsc_vld_n_outer_product_inst_bud),
      .out_product_rsc_rdy(out_product_rsc_rdy_n_tensor_weight_y_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn)
    );
  OpticalFlow_tensor_weight_y tensor_weight_y_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .out_product_rsc_dat(out_product_rsc_dat_n_outer_product_inst),
      .out_product_rsc_vld(out_product_rsc_vld_n_outer_product_inst_bud),
      .out_product_rsc_rdy(out_product_rsc_rdy_n_tensor_weight_y_inst_bud),
      .tensor_y_rsc_dat(tensor_y_rsc_dat_n_tensor_weight_y_inst),
      .tensor_y_rsc_vld(tensor_y_rsc_vld_n_tensor_weight_y_inst_bud),
      .tensor_y_rsc_rdy(tensor_y_rsc_rdy_n_tensor_weight_x_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .line_buf1_rsc_clken(line_buf1_rsc_clken_n_tensor_weight_y_inst),
      .line_buf1_rsc_q(line_buf1_rsc_tensor_weight_y_inst_q),
      .line_buf1_rsc_we(line_buf1_rsc_we_n_tensor_weight_y_inst_bud),
      .line_buf1_rsc_d(line_buf1_rsc_d_n_tensor_weight_y_inst),
      .line_buf1_rsc_adr(line_buf1_rsc_adr_n_tensor_weight_y_inst),
      .line_buf0_rsc_clken(line_buf0_rsc_clken_n_tensor_weight_y_inst),
      .line_buf0_rsc_q(line_buf0_rsc_tensor_weight_y_inst_q),
      .line_buf0_rsc_we(line_buf0_rsc_we_n_tensor_weight_y_inst_bud),
      .line_buf0_rsc_d(line_buf0_rsc_d_n_tensor_weight_y_inst),
      .line_buf0_rsc_adr(line_buf0_rsc_adr_n_tensor_weight_y_inst)
    );
  OpticalFlow_tensor_weight_x tensor_weight_x_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_y_rsc_dat(tensor_y_rsc_dat_n_tensor_weight_y_inst),
      .tensor_y_rsc_vld(tensor_y_rsc_vld_n_tensor_weight_y_inst_bud),
      .tensor_y_rsc_rdy(tensor_y_rsc_rdy_n_tensor_weight_x_inst_bud),
      .tensor_shift_rsc_dat(tensor_shift_rsc_dat_n_tensor_weight_x_inst),
      .tensor_shift_rsc_vld(tensor_shift_rsc_vld_n_tensor_weight_x_inst_bud),
      .tensor_shift_rsc_rdy(tensor_shift_rsc_rdy_n_flow_calc_inst_bud),
      .shift_rsc_dat(shift_rsc_dat_n_tensor_weight_x_inst),
      .shift_rsc_vld(shift_rsc_vld_n_tensor_weight_x_inst_bud),
      .shift_rsc_rdy(shift_rsc_rdy_n_flow_calc_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn)
    );
  OpticalFlow_flow_calc flow_calc_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .tensor_shift_rsc_dat(tensor_shift_rsc_dat_n_tensor_weight_x_inst),
      .tensor_shift_rsc_vld(tensor_shift_rsc_vld_n_tensor_weight_x_inst_bud),
      .tensor_shift_rsc_rdy(tensor_shift_rsc_rdy_n_flow_calc_inst_bud),
      .shift_rsc_dat(shift_rsc_dat_n_tensor_weight_x_inst),
      .shift_rsc_vld(shift_rsc_vld_n_tensor_weight_x_inst_bud),
      .shift_rsc_rdy(shift_rsc_rdy_n_flow_calc_inst_bud),
      .output_rsc_dat(output_rsc_dat_n_flow_calc_inst),
      .output_rsc_vld(output_rsc_vld_n_flow_calc_inst_bud),
      .output_rsc_rdy(outputs_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .shift_threshold(shift_threshold)
    );
  assign input_frames_rsc_rdy = input_frames_rsc_rdy_n_gradient_y_calc_inst_bud;
  assign line_buf3_rsc_clken = line_buf3_rsc_clken_n_gradient_y_calc_inst;
  assign line_buf3_rsc_we = line_buf3_rsc_we_n_gradient_y_calc_inst_bud;
  assign line_buf3_rsc_d = line_buf3_rsc_d_n_gradient_y_calc_inst;
  assign line_buf3_rsc_adr = line_buf3_rsc_adr_n_gradient_y_calc_inst;
  assign line_buf2_rsc_clken = line_buf2_rsc_clken_n_gradient_y_calc_inst;
  assign line_buf2_rsc_we = line_buf2_rsc_we_n_gradient_y_calc_inst_bud;
  assign line_buf2_rsc_d = line_buf2_rsc_d_n_gradient_y_calc_inst;
  assign line_buf2_rsc_adr = line_buf2_rsc_adr_n_gradient_y_calc_inst;
  assign line_buf1_rsc_gradient_y_calc_inst_clken = line_buf1_rsc_clken_n_gradient_y_calc_inst;
  assign line_buf1_rsc_gradient_y_calc_inst_we = line_buf1_rsc_we_n_gradient_y_calc_inst_bud;
  assign line_buf1_rsc_gradient_y_calc_inst_d = line_buf1_rsc_d_n_gradient_y_calc_inst;
  assign line_buf1_rsc_gradient_y_calc_inst_adr = line_buf1_rsc_adr_n_gradient_y_calc_inst;
  assign line_buf0_rsc_gradient_y_calc_inst_clken = line_buf0_rsc_clken_n_gradient_y_calc_inst;
  assign line_buf0_rsc_gradient_y_calc_inst_we = line_buf0_rsc_we_n_gradient_y_calc_inst_bud;
  assign line_buf0_rsc_gradient_y_calc_inst_d = line_buf0_rsc_d_n_gradient_y_calc_inst;
  assign line_buf0_rsc_gradient_y_calc_inst_adr = line_buf0_rsc_adr_n_gradient_y_calc_inst;
  assign line_buf5_Ix_rsc_clken = line_buf5_Ix_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf5_Ix_rsc_we = line_buf5_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf5_Ix_rsc_d = line_buf5_Ix_rsc_d_n_gradient_weight_y_inst;
  assign line_buf5_Ix_rsc_adr = line_buf5_Ix_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf4_Ix_rsc_clken = line_buf4_Ix_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf4_Ix_rsc_we = line_buf4_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf4_Ix_rsc_d = line_buf4_Ix_rsc_d_n_gradient_weight_y_inst;
  assign line_buf4_Ix_rsc_adr = line_buf4_Ix_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf3_Ix_rsc_clken = line_buf3_Ix_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf3_Ix_rsc_we = line_buf3_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf3_Ix_rsc_d = line_buf3_Ix_rsc_d_n_gradient_weight_y_inst;
  assign line_buf3_Ix_rsc_adr = line_buf3_Ix_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf2_Ix_rsc_clken = line_buf2_Ix_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf2_Ix_rsc_we = line_buf2_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf2_Ix_rsc_d = line_buf2_Ix_rsc_d_n_gradient_weight_y_inst;
  assign line_buf2_Ix_rsc_adr = line_buf2_Ix_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf1_Ix_rsc_clken = line_buf1_Ix_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf1_Ix_rsc_we = line_buf1_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf1_Ix_rsc_d = line_buf1_Ix_rsc_d_n_gradient_weight_y_inst;
  assign line_buf1_Ix_rsc_adr = line_buf1_Ix_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf0_Ix_rsc_clken = line_buf0_Ix_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf0_Ix_rsc_we = line_buf0_Ix_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf0_Ix_rsc_d = line_buf0_Ix_rsc_d_n_gradient_weight_y_inst;
  assign line_buf0_Ix_rsc_adr = line_buf0_Ix_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf5_Iy_rsc_clken = line_buf5_Iy_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf5_Iy_rsc_we = line_buf5_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf5_Iy_rsc_d = line_buf5_Iy_rsc_d_n_gradient_weight_y_inst;
  assign line_buf5_Iy_rsc_adr = line_buf5_Iy_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf4_Iy_rsc_clken = line_buf4_Iy_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf4_Iy_rsc_we = line_buf4_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf4_Iy_rsc_d = line_buf4_Iy_rsc_d_n_gradient_weight_y_inst;
  assign line_buf4_Iy_rsc_adr = line_buf4_Iy_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf3_Iy_rsc_clken = line_buf3_Iy_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf3_Iy_rsc_we = line_buf3_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf3_Iy_rsc_d = line_buf3_Iy_rsc_d_n_gradient_weight_y_inst;
  assign line_buf3_Iy_rsc_adr = line_buf3_Iy_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf2_Iy_rsc_clken = line_buf2_Iy_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf2_Iy_rsc_we = line_buf2_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf2_Iy_rsc_d = line_buf2_Iy_rsc_d_n_gradient_weight_y_inst;
  assign line_buf2_Iy_rsc_adr = line_buf2_Iy_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf1_Iy_rsc_clken = line_buf1_Iy_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf1_Iy_rsc_we = line_buf1_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf1_Iy_rsc_d = line_buf1_Iy_rsc_d_n_gradient_weight_y_inst;
  assign line_buf1_Iy_rsc_adr = line_buf1_Iy_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf0_Iy_rsc_clken = line_buf0_Iy_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf0_Iy_rsc_we = line_buf0_Iy_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf0_Iy_rsc_d = line_buf0_Iy_rsc_d_n_gradient_weight_y_inst;
  assign line_buf0_Iy_rsc_adr = line_buf0_Iy_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf5_Iz_rsc_clken = line_buf5_Iz_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf5_Iz_rsc_we = line_buf5_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf5_Iz_rsc_d = line_buf5_Iz_rsc_d_n_gradient_weight_y_inst;
  assign line_buf5_Iz_rsc_adr = line_buf5_Iz_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf4_Iz_rsc_clken = line_buf4_Iz_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf4_Iz_rsc_we = line_buf4_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf4_Iz_rsc_d = line_buf4_Iz_rsc_d_n_gradient_weight_y_inst;
  assign line_buf4_Iz_rsc_adr = line_buf4_Iz_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf3_Iz_rsc_clken = line_buf3_Iz_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf3_Iz_rsc_we = line_buf3_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf3_Iz_rsc_d = line_buf3_Iz_rsc_d_n_gradient_weight_y_inst;
  assign line_buf3_Iz_rsc_adr = line_buf3_Iz_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf2_Iz_rsc_clken = line_buf2_Iz_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf2_Iz_rsc_we = line_buf2_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf2_Iz_rsc_d = line_buf2_Iz_rsc_d_n_gradient_weight_y_inst;
  assign line_buf2_Iz_rsc_adr = line_buf2_Iz_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf1_Iz_rsc_clken = line_buf1_Iz_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf1_Iz_rsc_we = line_buf1_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf1_Iz_rsc_d = line_buf1_Iz_rsc_d_n_gradient_weight_y_inst;
  assign line_buf1_Iz_rsc_adr = line_buf1_Iz_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf0_Iz_rsc_clken = line_buf0_Iz_rsc_clken_n_gradient_weight_y_inst;
  assign line_buf0_Iz_rsc_we = line_buf0_Iz_rsc_we_n_gradient_weight_y_inst_bud;
  assign line_buf0_Iz_rsc_d = line_buf0_Iz_rsc_d_n_gradient_weight_y_inst;
  assign line_buf0_Iz_rsc_adr = line_buf0_Iz_rsc_adr_n_gradient_weight_y_inst;
  assign line_buf1_rsc_tensor_weight_y_inst_clken = line_buf1_rsc_clken_n_tensor_weight_y_inst;
  assign line_buf1_rsc_tensor_weight_y_inst_we = line_buf1_rsc_we_n_tensor_weight_y_inst_bud;
  assign line_buf1_rsc_tensor_weight_y_inst_d = line_buf1_rsc_d_n_tensor_weight_y_inst;
  assign line_buf1_rsc_tensor_weight_y_inst_adr = line_buf1_rsc_adr_n_tensor_weight_y_inst;
  assign line_buf0_rsc_tensor_weight_y_inst_clken = line_buf0_rsc_clken_n_tensor_weight_y_inst;
  assign line_buf0_rsc_tensor_weight_y_inst_we = line_buf0_rsc_we_n_tensor_weight_y_inst_bud;
  assign line_buf0_rsc_tensor_weight_y_inst_d = line_buf0_rsc_d_n_tensor_weight_y_inst;
  assign line_buf0_rsc_tensor_weight_y_inst_adr = line_buf0_rsc_adr_n_tensor_weight_y_inst;
  assign outputs_rsc_vld = output_rsc_vld_n_flow_calc_inst_bud;
  assign outputs_rsc_dat = output_rsc_dat_n_flow_calc_inst;
endmodule



